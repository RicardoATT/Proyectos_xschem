magic
tech sky130B
magscale 1 2
timestamp 1727994832
<< pwell >>
rect -2196 -279 2196 279
<< nmos >>
rect -2000 -131 2000 69
<< ndiff >>
rect -2058 57 -2000 69
rect -2058 -119 -2046 57
rect -2012 -119 -2000 57
rect -2058 -131 -2000 -119
rect 2000 57 2058 69
rect 2000 -119 2012 57
rect 2046 -119 2058 57
rect 2000 -131 2058 -119
<< ndiffc >>
rect -2046 -119 -2012 57
rect 2012 -119 2046 57
<< psubdiff >>
rect -2160 209 -2064 243
rect 2064 209 2160 243
rect -2160 147 -2126 209
rect 2126 147 2160 209
rect -2160 -209 -2126 -147
rect 2126 -209 2160 -147
rect -2160 -243 -2064 -209
rect 2064 -243 2160 -209
<< psubdiffcont >>
rect -2064 209 2064 243
rect -2160 -147 -2126 147
rect 2126 -147 2160 147
rect -2064 -243 2064 -209
<< poly >>
rect -2000 141 2000 157
rect -2000 107 -1984 141
rect 1984 107 2000 141
rect -2000 69 2000 107
rect -2000 -157 2000 -131
<< polycont >>
rect -1984 107 1984 141
<< locali >>
rect -2160 209 -2064 243
rect 2064 209 2160 243
rect -2160 147 -2126 209
rect 2126 147 2160 209
rect -2000 107 -1984 141
rect 1984 107 2000 141
rect -2046 57 -2012 73
rect -2046 -135 -2012 -119
rect 2012 57 2046 73
rect 2012 -135 2046 -119
rect -2160 -209 -2126 -147
rect 2126 -209 2160 -147
rect -2160 -243 -2064 -209
rect 2064 -243 2160 -209
<< viali >>
rect -1984 107 1984 141
rect -2046 -119 -2012 57
rect 2012 -119 2046 57
<< metal1 >>
rect -1996 141 1996 147
rect -1996 107 -1984 141
rect 1984 107 1996 141
rect -1996 101 1996 107
rect -2052 57 -2006 69
rect -2052 -119 -2046 57
rect -2012 -119 -2006 57
rect -2052 -131 -2006 -119
rect 2006 57 2052 69
rect 2006 -119 2012 57
rect 2046 -119 2052 57
rect 2006 -131 2052 -119
<< labels >>
flabel metal1 s -2029 -31 -2029 -31 0 FreeSans 480 0 0 0 D
port 0 nsew
flabel metal1 s -3 124 -3 124 0 FreeSans 480 0 0 0 G
port 1 nsew
flabel metal1 s 2029 -31 2029 -31 0 FreeSans 480 0 0 0 S
port 2 nsew
flabel locali s 2143 1 2143 1 0 FreeSans 480 0 0 0 B
port 3 nsew
<< properties >>
string FIXED_BBOX -2143 -226 2143 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 20.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
