magic
tech sky130B
magscale 1 2
timestamp 1728409957
<< error_s >>
rect 1268 1005 1303 1022
rect 1269 1004 1303 1005
rect 1269 968 1339 1004
rect 2625 968 2678 969
rect 1286 934 1357 968
rect 2607 934 2678 968
rect 1286 583 1356 934
rect 2608 933 2678 934
rect 2625 899 2696 933
rect 2976 899 3011 916
rect 1286 547 1339 583
rect 2625 530 2695 899
rect 2977 898 3011 899
rect 2977 862 3047 898
rect 2807 831 2865 837
rect 2807 797 2819 831
rect 2994 828 3065 862
rect 3345 828 3380 862
rect 2807 791 2865 797
rect 2807 613 2865 619
rect 2807 579 2819 613
rect 2807 573 2865 579
rect 2625 494 2678 530
rect 2994 477 3064 828
rect 3346 809 3380 828
rect 3176 760 3234 766
rect 3176 726 3188 760
rect 3176 720 3234 726
rect 3176 560 3234 566
rect 3176 526 3188 560
rect 3176 520 3234 526
rect 2994 441 3047 477
rect 3365 424 3380 809
rect 3399 775 3434 809
rect 3399 424 3433 775
rect 3545 707 3603 713
rect 3545 673 3557 707
rect 3545 667 3603 673
rect 3545 507 3603 513
rect 3545 473 3557 507
rect 3545 467 3603 473
rect 3399 390 3414 424
use sky130_fd_pr__pfet_01v8_HM8GCW  XM1
timestamp 1728409957
transform 1 0 643 0 1 811
box -696 -264 696 264
use sky130_fd_pr__nfet_01v8_43PFCA  XM2
timestamp 1728409957
transform 1 0 1982 0 1 749
box -696 -255 696 255
use sky130_fd_pr__pfet_01v8_MJH8BZ  XM3
timestamp 1728409957
transform 1 0 2836 0 1 705
box -211 -264 211 264
use sky130_fd_pr__nfet_01v8_HVW3BE  XM4
timestamp 1728409957
transform 1 0 3205 0 1 643
box -211 -255 211 255
use sky130_fd_pr__nfet_01v8_HVW3BE  XM5
timestamp 1728409957
transform 1 0 3574 0 1 590
box -211 -255 211 255
<< end >>
