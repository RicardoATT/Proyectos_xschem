magic
tech sky130B
magscale 1 2
timestamp 1728434276
<< error_p >>
rect -29 1572 29 1578
rect -29 1538 -17 1572
rect -29 1532 29 1538
rect -29 -1538 29 -1532
rect -29 -1572 -17 -1538
rect -29 -1578 29 -1572
<< pwell >>
rect -211 -1710 211 1710
<< nmos >>
rect -15 -1500 15 1500
<< ndiff >>
rect -73 1488 -15 1500
rect -73 -1488 -61 1488
rect -27 -1488 -15 1488
rect -73 -1500 -15 -1488
rect 15 1488 73 1500
rect 15 -1488 27 1488
rect 61 -1488 73 1488
rect 15 -1500 73 -1488
<< ndiffc >>
rect -61 -1488 -27 1488
rect 27 -1488 61 1488
<< psubdiff >>
rect -175 1640 -79 1674
rect 79 1640 175 1674
rect -175 1578 -141 1640
rect 141 1578 175 1640
rect -175 -1640 -141 -1578
rect 141 -1640 175 -1578
rect -175 -1674 -79 -1640
rect 79 -1674 175 -1640
<< psubdiffcont >>
rect -79 1640 79 1674
rect -175 -1578 -141 1578
rect 141 -1578 175 1578
rect -79 -1674 79 -1640
<< poly >>
rect -33 1572 33 1588
rect -33 1538 -17 1572
rect 17 1538 33 1572
rect -33 1522 33 1538
rect -15 1500 15 1522
rect -15 -1522 15 -1500
rect -33 -1538 33 -1522
rect -33 -1572 -17 -1538
rect 17 -1572 33 -1538
rect -33 -1588 33 -1572
<< polycont >>
rect -17 1538 17 1572
rect -17 -1572 17 -1538
<< locali >>
rect -175 1640 -79 1674
rect 79 1640 175 1674
rect -175 1578 -141 1640
rect 141 1578 175 1640
rect -33 1538 -17 1572
rect 17 1538 33 1572
rect -61 1488 -27 1504
rect -61 -1504 -27 -1488
rect 27 1488 61 1504
rect 27 -1504 61 -1488
rect -33 -1572 -17 -1538
rect 17 -1572 33 -1538
rect -175 -1640 -141 -1578
rect 141 -1640 175 -1578
rect -175 -1674 -79 -1640
rect 79 -1674 175 -1640
<< viali >>
rect -17 1538 17 1572
rect -61 -1488 -27 1488
rect 27 -1488 61 1488
rect -17 -1572 17 -1538
<< metal1 >>
rect -29 1572 29 1578
rect -29 1538 -17 1572
rect 17 1538 29 1572
rect -29 1532 29 1538
rect -67 1488 -21 1500
rect -67 -1488 -61 1488
rect -27 -1488 -21 1488
rect -67 -1500 -21 -1488
rect 21 1488 67 1500
rect 21 -1488 27 1488
rect 61 -1488 67 1488
rect 21 -1500 67 -1488
rect -29 -1538 29 -1532
rect -29 -1572 -17 -1538
rect 17 -1572 29 -1538
rect -29 -1578 29 -1572
<< properties >>
string FIXED_BBOX -158 -1657 158 1657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 15.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
