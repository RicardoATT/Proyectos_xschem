magic
tech sky130B
magscale 1 2
timestamp 1728522838
<< locali >>
rect 555 8589 623 9785
rect 23 8475 101 8509
rect 355 8273 389 8307
rect -7 8201 27 8273
rect 355 8167 389 8201
rect 575 8089 609 8182
rect 12 8053 101 8087
rect 418 6881 495 6915
rect -7 6103 27 6213
rect 485 6166 519 6276
rect 379 6103 413 6137
rect 485 6103 490 6137
rect 485 5491 519 5611
rect 757 5407 791 5484
rect 299 4959 379 4993
rect -7 4691 27 4811
rect -7 4159 27 4245
rect 485 4138 519 4258
rect 195 3600 229 3690
rect -7 3537 61 3578
rect 339 3573 579 3607
rect 617 3604 651 3696
rect 731 3573 4432 3607
<< viali >>
rect 384 6881 418 6915
rect 4432 3573 4466 3607
<< metal1 >>
rect 492 8433 541 8477
rect 371 8307 405 8421
rect 489 8419 541 8433
rect 507 8369 541 8419
rect 492 8317 498 8369
rect 550 8317 556 8369
rect 371 8273 462 8307
rect 346 8210 398 8216
rect 346 8152 398 8158
rect 252 7073 286 7090
rect 233 7045 286 7073
rect 67 6989 117 7029
rect -16 6804 36 6810
rect -16 6746 36 6752
rect -7 6209 27 6746
rect 67 6593 101 6989
rect 233 6693 267 7045
rect 355 6983 389 8152
rect 428 7019 462 8273
rect 507 8216 541 8317
rect 498 8210 550 8216
rect 498 8152 550 8158
rect 309 6955 389 6983
rect 419 7013 471 7019
rect 419 6955 471 6961
rect 309 6810 343 6955
rect 378 6915 424 6927
rect 378 6881 384 6915
rect 418 6881 424 6915
rect 378 6869 424 6881
rect 300 6804 352 6810
rect 300 6746 352 6752
rect 185 6659 267 6693
rect 107 6041 141 6363
rect 195 6137 229 6354
rect 386 6219 415 6869
rect 368 6167 374 6219
rect 426 6167 432 6219
rect 195 6103 369 6137
rect 107 6001 169 6041
rect 335 5405 369 6103
rect 507 5725 541 8152
rect 663 7089 835 7117
rect 643 6697 677 7042
rect 801 6659 835 7089
rect 721 6631 835 6659
rect 599 6190 633 6413
rect 678 6305 730 6311
rect 678 6247 730 6253
rect 590 6184 642 6190
rect 590 6126 642 6132
rect 599 6058 633 6126
rect 687 6055 721 6247
rect 507 5691 650 5725
rect 801 5623 835 6631
rect 801 5589 4484 5623
rect 801 5517 835 5589
rect 801 5483 905 5517
rect 335 5377 593 5405
rect 373 5330 425 5336
rect 373 5272 425 5278
rect 492 5275 498 5327
rect 550 5275 556 5327
rect -16 4934 36 4940
rect -43 4891 -16 4925
rect 204 4891 343 4925
rect -16 4876 36 4882
rect 177 4832 229 4838
rect -43 4789 177 4823
rect 177 4774 229 4780
rect 94 4726 154 4739
rect 94 4674 98 4726
rect 150 4717 154 4726
rect 309 4717 343 4891
rect 150 4683 343 4717
rect 150 4674 154 4683
rect 94 4661 154 4674
rect 107 4605 141 4661
rect 384 4605 413 5272
rect 229 4576 413 4605
rect 300 4522 352 4528
rect 300 4464 352 4470
rect -43 4333 185 4367
rect 309 4274 343 4464
rect 309 4222 370 4274
rect 422 4222 428 4274
rect 507 4159 541 5275
rect 678 4274 712 4367
rect 663 4222 669 4274
rect 721 4222 727 4274
rect -43 4125 27 4159
rect -7 4057 27 4125
rect 415 4125 541 4159
rect -7 4023 197 4057
rect 415 3985 449 4125
rect 871 4057 905 5483
rect 604 4023 905 4057
rect 101 3957 141 3985
rect 415 3951 563 3985
rect -16 3725 36 3731
rect 36 3685 102 3713
rect -16 3667 36 3673
rect 4419 3616 4479 3629
rect 4419 3564 4423 3616
rect 4475 3564 4479 3616
rect 4419 3551 4479 3564
<< via1 >>
rect 498 8317 550 8369
rect 346 8158 398 8210
rect -16 6752 36 6804
rect 498 8158 550 8210
rect 419 6961 471 7013
rect 300 6752 352 6804
rect 374 6167 426 6219
rect 678 6253 730 6305
rect 590 6132 642 6184
rect 373 5278 425 5330
rect 498 5275 550 5327
rect -16 4882 36 4934
rect 177 4780 229 4832
rect 98 4674 150 4726
rect 300 4470 352 4522
rect 370 4222 422 4274
rect 669 4222 721 4274
rect -16 3673 36 3725
rect 4423 3607 4475 3616
rect 4423 3573 4432 3607
rect 4432 3573 4466 3607
rect 4466 3573 4475 3607
rect 4423 3564 4475 3573
<< metal2 >>
rect 29 8313 38 8373
rect 98 8360 107 8373
rect 498 8369 550 8375
rect 98 8326 498 8360
rect 98 8313 107 8326
rect 498 8311 550 8317
rect 340 8158 346 8210
rect 398 8201 404 8210
rect 492 8201 498 8210
rect 398 8167 498 8201
rect 398 8158 404 8167
rect 492 8158 498 8167
rect 550 8158 556 8210
rect 419 7013 471 7019
rect 419 6955 471 6961
rect -22 6752 -16 6804
rect 36 6795 42 6804
rect 294 6795 300 6804
rect 36 6761 300 6795
rect 36 6752 42 6761
rect 294 6752 300 6761
rect 352 6752 358 6804
rect 428 6296 462 6955
rect 672 6296 678 6305
rect 428 6262 678 6296
rect 672 6253 678 6262
rect 730 6253 736 6305
rect 374 6219 426 6225
rect 584 6175 590 6184
rect 374 6161 426 6167
rect 385 5330 414 6161
rect 507 6141 590 6175
rect 507 5333 541 6141
rect 584 6132 590 6141
rect 642 6132 648 6184
rect 367 5278 373 5330
rect 425 5278 431 5330
rect 498 5327 550 5333
rect 498 5269 550 5275
rect -22 4882 -16 4934
rect 36 4882 42 4934
rect -7 3731 27 4882
rect 171 4780 177 4832
rect 229 4823 235 4832
rect 229 4789 343 4823
rect 229 4780 235 4789
rect 94 4730 154 4739
rect 94 4661 154 4670
rect 309 4522 343 4789
rect 294 4470 300 4522
rect 352 4470 358 4522
rect 669 4274 721 4280
rect 364 4222 370 4274
rect 422 4265 428 4274
rect 422 4231 669 4265
rect 422 4222 428 4231
rect 669 4216 721 4222
rect -16 3725 36 3731
rect -16 3667 36 3673
rect 4419 3620 4479 3629
rect 4419 3551 4479 3560
<< via2 >>
rect 38 8313 98 8373
rect 94 4726 154 4730
rect 94 4674 98 4726
rect 98 4674 150 4726
rect 150 4674 154 4726
rect 94 4670 154 4674
rect 4419 3616 4479 3620
rect 4419 3564 4423 3616
rect 4423 3564 4475 3616
rect 4475 3564 4479 3616
rect 4419 3560 4479 3564
<< metal3 >>
rect 33 8373 103 8378
rect 33 8313 38 8373
rect 98 8313 103 8373
rect 33 8308 103 8313
rect 38 8167 98 8308
rect 89 4730 159 4735
rect 89 4670 94 4730
rect 154 4670 246 4730
rect 89 4665 159 4670
rect 4417 3788 4481 3794
rect 4417 3718 4481 3724
rect 4419 3625 4479 3718
rect 4414 3620 4484 3625
rect 4414 3560 4419 3620
rect 4479 3560 4484 3620
rect 4414 3555 4484 3560
<< via3 >>
rect 4417 3724 4481 3788
<< metal4 >>
rect 4167 5516 4227 5892
rect 4416 3788 4482 3789
rect 4416 3786 4417 3788
rect 4167 3726 4417 3786
rect 4416 3724 4417 3726
rect 4481 3724 4482 3788
rect 4416 3723 4482 3724
use sky130_fd_pr__cap_mim_m3_1_BNHTNG  sky130_fd_pr__cap_mim_m3_1_BNHTNG_0
timestamp 1728522838
transform -1 0 2143 0 1 7745
box -2186 -2040 2186 2040
use sky130_fd_pr__cap_mim_m3_1_TNHPNJ  sky130_fd_pr__cap_mim_m3_1_TNHPNJ_0
timestamp 1728522838
transform -1 0 2143 0 1 4577
box -2186 -1040 2186 1040
use sky130_fd_pr__nfet_01v8_8TTSKH  sky130_fd_pr__nfet_01v8_8TTSKH_0
timestamp 1728500067
transform 1 0 695 0 -1 4874
box -246 -679 246 679
use sky130_fd_pr__nfet_01v8_84Z3BM  sky130_fd_pr__nfet_01v8_84Z3BM_0
timestamp 1728500067
transform -1 0 660 0 1 6540
box -211 -329 211 329
use sky130_fd_pr__nfet_01v8_84Z3BM  XM1
timestamp 1728500067
transform 1 0 168 0 1 3866
box -211 -329 211 329
use sky130_fd_pr__nfet_01v8_8TEW3F  XM2
timestamp 1728522838
transform 1 0 203 0 1 5463
box -246 -710 246 710
use sky130_fd_pr__pfet_01v8_FQSSVM  XM3
timestamp 1728501028
transform 0 -1 191 1 0 7541
box -696 -234 696 234
use sky130_fd_pr__nfet_01v8_84Z3BM  XM4
timestamp 1728500067
transform 1 0 168 0 1 6502
box -211 -329 211 329
use sky130_fd_pr__pfet_01v8_LJP3BL  XM6
timestamp 1728501028
transform 0 -1 291 1 0 8448
box -211 -334 211 334
use sky130_fd_pr__nfet_01v8_84Z3BM  XM7
timestamp 1728500067
transform -1 0 660 0 -1 5882
box -211 -329 211 329
use sky130_fd_pr__pfet_01v8_MGSVTG  XM8
timestamp 1728501028
transform -1 0 636 0 1 7553
box -211 -684 211 684
use sky130_fd_pr__nfet_01v8_84Z3BM  XM10
timestamp 1728500067
transform 1 0 590 0 1 3866
box -211 -329 211 329
use sky130_fd_pr__nfet_01v8_64Z3AY  XM11
timestamp 1728500067
transform -1 0 168 0 -1 4474
box -211 -279 211 279
<< labels >>
flabel metal1 s -43 4789 -43 4823 0 FreeSans 480 0 0 0 Vb
port 2 nsew
flabel metal1 s -43 4891 -43 4925 0 FreeSans 480 0 0 0 Iin
port 3 nsew
flabel metal1 s -43 4333 -43 4367 0 FreeSans 480 0 0 0 Vinh
port 4 nsew
flabel metal1 s -43 4125 -43 4159 0 FreeSans 480 0 0 0 Vlky
port 5 nsew
flabel locali s 555 9785 623 9785 0 FreeSans 480 0 0 0 VDD
port 8 nsew
flabel locali s -7 3537 61 3537 0 FreeSans 480 0 0 0 GND
port 9 nsew
flabel metal1 s 4484 5589 4484 5623 0 FreeSans 480 0 0 0 Vout
port 10 nsew
<< end >>
