*MADE BY JORGE ALEJANDRO JUAREZ LORA IPN

.subckt rram_v1 TE BE
N1 TE BE rram_v1_model gap_initial=unif(0.9,0.8)
.ends rram_v1

.model rram_v1_model rram_v1_va


.control
pre_osdi /home/ricardo/pdk/sky130B/libs.tech/ngspice/rram_v1.osdi
.endc
