magic
tech sky130B
magscale 1 2
timestamp 1729119800
<< error_p >>
rect -845 231 -787 237
rect -653 231 -595 237
rect -461 231 -403 237
rect -269 231 -211 237
rect -77 231 -19 237
rect 115 231 173 237
rect 307 231 365 237
rect 499 231 557 237
rect 691 231 749 237
rect 883 231 941 237
rect -845 197 -833 231
rect -653 197 -641 231
rect -461 197 -449 231
rect -269 197 -257 231
rect -77 197 -65 231
rect 115 197 127 231
rect 307 197 319 231
rect 499 197 511 231
rect 691 197 703 231
rect 883 197 895 231
rect -845 191 -787 197
rect -653 191 -595 197
rect -461 191 -403 197
rect -269 191 -211 197
rect -77 191 -19 197
rect 115 191 173 197
rect 307 191 365 197
rect 499 191 557 197
rect 691 191 749 197
rect 883 191 941 197
rect -941 -197 -883 -191
rect -749 -197 -691 -191
rect -557 -197 -499 -191
rect -365 -197 -307 -191
rect -173 -197 -115 -191
rect 19 -197 77 -191
rect 211 -197 269 -191
rect 403 -197 461 -191
rect 595 -197 653 -191
rect 787 -197 845 -191
rect -941 -231 -929 -197
rect -749 -231 -737 -197
rect -557 -231 -545 -197
rect -365 -231 -353 -197
rect -173 -231 -161 -197
rect 19 -231 31 -197
rect 211 -231 223 -197
rect 403 -231 415 -197
rect 595 -231 607 -197
rect 787 -231 799 -197
rect -941 -237 -883 -231
rect -749 -237 -691 -231
rect -557 -237 -499 -231
rect -365 -237 -307 -231
rect -173 -237 -115 -231
rect 19 -237 77 -231
rect 211 -237 269 -231
rect 403 -237 461 -231
rect 595 -237 653 -231
rect 787 -237 845 -231
<< nwell >>
rect -1127 -369 1127 369
<< pmos >>
rect -927 -150 -897 150
rect -831 -150 -801 150
rect -735 -150 -705 150
rect -639 -150 -609 150
rect -543 -150 -513 150
rect -447 -150 -417 150
rect -351 -150 -321 150
rect -255 -150 -225 150
rect -159 -150 -129 150
rect -63 -150 -33 150
rect 33 -150 63 150
rect 129 -150 159 150
rect 225 -150 255 150
rect 321 -150 351 150
rect 417 -150 447 150
rect 513 -150 543 150
rect 609 -150 639 150
rect 705 -150 735 150
rect 801 -150 831 150
rect 897 -150 927 150
<< pdiff >>
rect -989 138 -927 150
rect -989 -138 -977 138
rect -943 -138 -927 138
rect -989 -150 -927 -138
rect -897 138 -831 150
rect -897 -138 -881 138
rect -847 -138 -831 138
rect -897 -150 -831 -138
rect -801 138 -735 150
rect -801 -138 -785 138
rect -751 -138 -735 138
rect -801 -150 -735 -138
rect -705 138 -639 150
rect -705 -138 -689 138
rect -655 -138 -639 138
rect -705 -150 -639 -138
rect -609 138 -543 150
rect -609 -138 -593 138
rect -559 -138 -543 138
rect -609 -150 -543 -138
rect -513 138 -447 150
rect -513 -138 -497 138
rect -463 -138 -447 138
rect -513 -150 -447 -138
rect -417 138 -351 150
rect -417 -138 -401 138
rect -367 -138 -351 138
rect -417 -150 -351 -138
rect -321 138 -255 150
rect -321 -138 -305 138
rect -271 -138 -255 138
rect -321 -150 -255 -138
rect -225 138 -159 150
rect -225 -138 -209 138
rect -175 -138 -159 138
rect -225 -150 -159 -138
rect -129 138 -63 150
rect -129 -138 -113 138
rect -79 -138 -63 138
rect -129 -150 -63 -138
rect -33 138 33 150
rect -33 -138 -17 138
rect 17 -138 33 138
rect -33 -150 33 -138
rect 63 138 129 150
rect 63 -138 79 138
rect 113 -138 129 138
rect 63 -150 129 -138
rect 159 138 225 150
rect 159 -138 175 138
rect 209 -138 225 138
rect 159 -150 225 -138
rect 255 138 321 150
rect 255 -138 271 138
rect 305 -138 321 138
rect 255 -150 321 -138
rect 351 138 417 150
rect 351 -138 367 138
rect 401 -138 417 138
rect 351 -150 417 -138
rect 447 138 513 150
rect 447 -138 463 138
rect 497 -138 513 138
rect 447 -150 513 -138
rect 543 138 609 150
rect 543 -138 559 138
rect 593 -138 609 138
rect 543 -150 609 -138
rect 639 138 705 150
rect 639 -138 655 138
rect 689 -138 705 138
rect 639 -150 705 -138
rect 735 138 801 150
rect 735 -138 751 138
rect 785 -138 801 138
rect 735 -150 801 -138
rect 831 138 897 150
rect 831 -138 847 138
rect 881 -138 897 138
rect 831 -150 897 -138
rect 927 138 989 150
rect 927 -138 943 138
rect 977 -138 989 138
rect 927 -150 989 -138
<< pdiffc >>
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
<< nsubdiff >>
rect -1091 299 -995 333
rect 995 299 1091 333
rect -1091 237 -1057 299
rect 1057 237 1091 299
rect -1091 -299 -1057 -237
rect 1057 -299 1091 -237
rect -1091 -333 -995 -299
rect 995 -333 1091 -299
<< nsubdiffcont >>
rect -995 299 995 333
rect -1091 -237 -1057 237
rect 1057 -237 1091 237
rect -995 -333 995 -299
<< poly >>
rect -849 231 -783 247
rect -849 197 -833 231
rect -799 197 -783 231
rect -849 181 -783 197
rect -657 231 -591 247
rect -657 197 -641 231
rect -607 197 -591 231
rect -657 181 -591 197
rect -465 231 -399 247
rect -465 197 -449 231
rect -415 197 -399 231
rect -465 181 -399 197
rect -273 231 -207 247
rect -273 197 -257 231
rect -223 197 -207 231
rect -273 181 -207 197
rect -81 231 -15 247
rect -81 197 -65 231
rect -31 197 -15 231
rect -81 181 -15 197
rect 111 231 177 247
rect 111 197 127 231
rect 161 197 177 231
rect 111 181 177 197
rect 303 231 369 247
rect 303 197 319 231
rect 353 197 369 231
rect 303 181 369 197
rect 495 231 561 247
rect 495 197 511 231
rect 545 197 561 231
rect 495 181 561 197
rect 687 231 753 247
rect 687 197 703 231
rect 737 197 753 231
rect 687 181 753 197
rect 879 231 945 247
rect 879 197 895 231
rect 929 197 945 231
rect 879 181 945 197
rect -927 150 -897 176
rect -831 150 -801 181
rect -735 150 -705 176
rect -639 150 -609 181
rect -543 150 -513 176
rect -447 150 -417 181
rect -351 150 -321 176
rect -255 150 -225 181
rect -159 150 -129 176
rect -63 150 -33 181
rect 33 150 63 176
rect 129 150 159 181
rect 225 150 255 176
rect 321 150 351 181
rect 417 150 447 176
rect 513 150 543 181
rect 609 150 639 176
rect 705 150 735 181
rect 801 150 831 176
rect 897 150 927 181
rect -927 -181 -897 -150
rect -831 -176 -801 -150
rect -735 -181 -705 -150
rect -639 -176 -609 -150
rect -543 -181 -513 -150
rect -447 -176 -417 -150
rect -351 -181 -321 -150
rect -255 -176 -225 -150
rect -159 -181 -129 -150
rect -63 -176 -33 -150
rect 33 -181 63 -150
rect 129 -176 159 -150
rect 225 -181 255 -150
rect 321 -176 351 -150
rect 417 -181 447 -150
rect 513 -176 543 -150
rect 609 -181 639 -150
rect 705 -176 735 -150
rect 801 -181 831 -150
rect 897 -176 927 -150
rect -945 -197 -879 -181
rect -945 -231 -929 -197
rect -895 -231 -879 -197
rect -945 -247 -879 -231
rect -753 -197 -687 -181
rect -753 -231 -737 -197
rect -703 -231 -687 -197
rect -753 -247 -687 -231
rect -561 -197 -495 -181
rect -561 -231 -545 -197
rect -511 -231 -495 -197
rect -561 -247 -495 -231
rect -369 -197 -303 -181
rect -369 -231 -353 -197
rect -319 -231 -303 -197
rect -369 -247 -303 -231
rect -177 -197 -111 -181
rect -177 -231 -161 -197
rect -127 -231 -111 -197
rect -177 -247 -111 -231
rect 15 -197 81 -181
rect 15 -231 31 -197
rect 65 -231 81 -197
rect 15 -247 81 -231
rect 207 -197 273 -181
rect 207 -231 223 -197
rect 257 -231 273 -197
rect 207 -247 273 -231
rect 399 -197 465 -181
rect 399 -231 415 -197
rect 449 -231 465 -197
rect 399 -247 465 -231
rect 591 -197 657 -181
rect 591 -231 607 -197
rect 641 -231 657 -197
rect 591 -247 657 -231
rect 783 -197 849 -181
rect 783 -231 799 -197
rect 833 -231 849 -197
rect 783 -247 849 -231
<< polycont >>
rect -833 197 -799 231
rect -641 197 -607 231
rect -449 197 -415 231
rect -257 197 -223 231
rect -65 197 -31 231
rect 127 197 161 231
rect 319 197 353 231
rect 511 197 545 231
rect 703 197 737 231
rect 895 197 929 231
rect -929 -231 -895 -197
rect -737 -231 -703 -197
rect -545 -231 -511 -197
rect -353 -231 -319 -197
rect -161 -231 -127 -197
rect 31 -231 65 -197
rect 223 -231 257 -197
rect 415 -231 449 -197
rect 607 -231 641 -197
rect 799 -231 833 -197
<< locali >>
rect -1091 299 -995 333
rect 995 299 1091 333
rect -1091 237 -1057 299
rect 1057 237 1091 299
rect -849 197 -833 231
rect -799 197 -783 231
rect -657 197 -641 231
rect -607 197 -591 231
rect -465 197 -449 231
rect -415 197 -399 231
rect -273 197 -257 231
rect -223 197 -207 231
rect -81 197 -65 231
rect -31 197 -15 231
rect 111 197 127 231
rect 161 197 177 231
rect 303 197 319 231
rect 353 197 369 231
rect 495 197 511 231
rect 545 197 561 231
rect 687 197 703 231
rect 737 197 753 231
rect 879 197 895 231
rect 929 197 945 231
rect -977 138 -943 154
rect -977 -154 -943 -138
rect -881 138 -847 154
rect -881 -154 -847 -138
rect -785 138 -751 154
rect -785 -154 -751 -138
rect -689 138 -655 154
rect -689 -154 -655 -138
rect -593 138 -559 154
rect -593 -154 -559 -138
rect -497 138 -463 154
rect -497 -154 -463 -138
rect -401 138 -367 154
rect -401 -154 -367 -138
rect -305 138 -271 154
rect -305 -154 -271 -138
rect -209 138 -175 154
rect -209 -154 -175 -138
rect -113 138 -79 154
rect -113 -154 -79 -138
rect -17 138 17 154
rect -17 -154 17 -138
rect 79 138 113 154
rect 79 -154 113 -138
rect 175 138 209 154
rect 175 -154 209 -138
rect 271 138 305 154
rect 271 -154 305 -138
rect 367 138 401 154
rect 367 -154 401 -138
rect 463 138 497 154
rect 463 -154 497 -138
rect 559 138 593 154
rect 559 -154 593 -138
rect 655 138 689 154
rect 655 -154 689 -138
rect 751 138 785 154
rect 751 -154 785 -138
rect 847 138 881 154
rect 847 -154 881 -138
rect 943 138 977 154
rect 943 -154 977 -138
rect -945 -231 -929 -197
rect -895 -231 -879 -197
rect -753 -231 -737 -197
rect -703 -231 -687 -197
rect -561 -231 -545 -197
rect -511 -231 -495 -197
rect -369 -231 -353 -197
rect -319 -231 -303 -197
rect -177 -231 -161 -197
rect -127 -231 -111 -197
rect 15 -231 31 -197
rect 65 -231 81 -197
rect 207 -231 223 -197
rect 257 -231 273 -197
rect 399 -231 415 -197
rect 449 -231 465 -197
rect 591 -231 607 -197
rect 641 -231 657 -197
rect 783 -231 799 -197
rect 833 -231 849 -197
rect -1091 -299 -1057 -237
rect 1057 -299 1091 -237
rect -1091 -333 -995 -299
rect 995 -333 1091 -299
<< viali >>
rect -833 197 -799 231
rect -641 197 -607 231
rect -449 197 -415 231
rect -257 197 -223 231
rect -65 197 -31 231
rect 127 197 161 231
rect 319 197 353 231
rect 511 197 545 231
rect 703 197 737 231
rect 895 197 929 231
rect -977 -138 -943 138
rect -881 -138 -847 138
rect -785 -138 -751 138
rect -689 -138 -655 138
rect -593 -138 -559 138
rect -497 -138 -463 138
rect -401 -138 -367 138
rect -305 -138 -271 138
rect -209 -138 -175 138
rect -113 -138 -79 138
rect -17 -138 17 138
rect 79 -138 113 138
rect 175 -138 209 138
rect 271 -138 305 138
rect 367 -138 401 138
rect 463 -138 497 138
rect 559 -138 593 138
rect 655 -138 689 138
rect 751 -138 785 138
rect 847 -138 881 138
rect 943 -138 977 138
rect -929 -231 -895 -197
rect -737 -231 -703 -197
rect -545 -231 -511 -197
rect -353 -231 -319 -197
rect -161 -231 -127 -197
rect 31 -231 65 -197
rect 223 -231 257 -197
rect 415 -231 449 -197
rect 607 -231 641 -197
rect 799 -231 833 -197
<< metal1 >>
rect -845 231 -787 237
rect -845 197 -833 231
rect -799 197 -787 231
rect -845 191 -787 197
rect -653 231 -595 237
rect -653 197 -641 231
rect -607 197 -595 231
rect -653 191 -595 197
rect -461 231 -403 237
rect -461 197 -449 231
rect -415 197 -403 231
rect -461 191 -403 197
rect -269 231 -211 237
rect -269 197 -257 231
rect -223 197 -211 231
rect -269 191 -211 197
rect -77 231 -19 237
rect -77 197 -65 231
rect -31 197 -19 231
rect -77 191 -19 197
rect 115 231 173 237
rect 115 197 127 231
rect 161 197 173 231
rect 115 191 173 197
rect 307 231 365 237
rect 307 197 319 231
rect 353 197 365 231
rect 307 191 365 197
rect 499 231 557 237
rect 499 197 511 231
rect 545 197 557 231
rect 499 191 557 197
rect 691 231 749 237
rect 691 197 703 231
rect 737 197 749 231
rect 691 191 749 197
rect 883 231 941 237
rect 883 197 895 231
rect 929 197 941 231
rect 883 191 941 197
rect -983 138 -937 150
rect -983 -138 -977 138
rect -943 -138 -937 138
rect -983 -150 -937 -138
rect -887 138 -841 150
rect -887 -138 -881 138
rect -847 -138 -841 138
rect -887 -150 -841 -138
rect -791 138 -745 150
rect -791 -138 -785 138
rect -751 -138 -745 138
rect -791 -150 -745 -138
rect -695 138 -649 150
rect -695 -138 -689 138
rect -655 -138 -649 138
rect -695 -150 -649 -138
rect -599 138 -553 150
rect -599 -138 -593 138
rect -559 -138 -553 138
rect -599 -150 -553 -138
rect -503 138 -457 150
rect -503 -138 -497 138
rect -463 -138 -457 138
rect -503 -150 -457 -138
rect -407 138 -361 150
rect -407 -138 -401 138
rect -367 -138 -361 138
rect -407 -150 -361 -138
rect -311 138 -265 150
rect -311 -138 -305 138
rect -271 -138 -265 138
rect -311 -150 -265 -138
rect -215 138 -169 150
rect -215 -138 -209 138
rect -175 -138 -169 138
rect -215 -150 -169 -138
rect -119 138 -73 150
rect -119 -138 -113 138
rect -79 -138 -73 138
rect -119 -150 -73 -138
rect -23 138 23 150
rect -23 -138 -17 138
rect 17 -138 23 138
rect -23 -150 23 -138
rect 73 138 119 150
rect 73 -138 79 138
rect 113 -138 119 138
rect 73 -150 119 -138
rect 169 138 215 150
rect 169 -138 175 138
rect 209 -138 215 138
rect 169 -150 215 -138
rect 265 138 311 150
rect 265 -138 271 138
rect 305 -138 311 138
rect 265 -150 311 -138
rect 361 138 407 150
rect 361 -138 367 138
rect 401 -138 407 138
rect 361 -150 407 -138
rect 457 138 503 150
rect 457 -138 463 138
rect 497 -138 503 138
rect 457 -150 503 -138
rect 553 138 599 150
rect 553 -138 559 138
rect 593 -138 599 138
rect 553 -150 599 -138
rect 649 138 695 150
rect 649 -138 655 138
rect 689 -138 695 138
rect 649 -150 695 -138
rect 745 138 791 150
rect 745 -138 751 138
rect 785 -138 791 138
rect 745 -150 791 -138
rect 841 138 887 150
rect 841 -138 847 138
rect 881 -138 887 138
rect 841 -150 887 -138
rect 937 138 983 150
rect 937 -138 943 138
rect 977 -138 983 138
rect 937 -150 983 -138
rect -941 -197 -883 -191
rect -941 -231 -929 -197
rect -895 -231 -883 -197
rect -941 -237 -883 -231
rect -749 -197 -691 -191
rect -749 -231 -737 -197
rect -703 -231 -691 -197
rect -749 -237 -691 -231
rect -557 -197 -499 -191
rect -557 -231 -545 -197
rect -511 -231 -499 -197
rect -557 -237 -499 -231
rect -365 -197 -307 -191
rect -365 -231 -353 -197
rect -319 -231 -307 -197
rect -365 -237 -307 -231
rect -173 -197 -115 -191
rect -173 -231 -161 -197
rect -127 -231 -115 -197
rect -173 -237 -115 -231
rect 19 -197 77 -191
rect 19 -231 31 -197
rect 65 -231 77 -197
rect 19 -237 77 -231
rect 211 -197 269 -191
rect 211 -231 223 -197
rect 257 -231 269 -197
rect 211 -237 269 -231
rect 403 -197 461 -191
rect 403 -231 415 -197
rect 449 -231 461 -197
rect 403 -237 461 -231
rect 595 -197 653 -191
rect 595 -231 607 -197
rect 641 -231 653 -197
rect 595 -237 653 -231
rect 787 -197 845 -191
rect 787 -231 799 -197
rect 833 -231 845 -197
rect 787 -237 845 -231
<< properties >>
string FIXED_BBOX -1074 -316 1074 316
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
