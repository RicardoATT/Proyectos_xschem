magic
tech sky130B
magscale 1 2
timestamp 1728608927
<< locali >>
rect 3563 8648 3633 8718
rect 3101 8534 3297 8568
rect 3597 7682 4125 7692
rect 3563 7658 4125 7682
rect 4091 7608 4125 7658
rect 4293 7503 4327 7642
rect 3669 6930 3703 7070
rect 3871 7036 3905 7160
rect 4091 6940 4125 7080
rect 4205 6825 4239 6974
rect 3669 6272 3703 6412
rect 3669 5614 3703 5754
rect 4091 4914 4125 5054
rect 2543 4326 2613 4396
rect 2651 4362 2687 4510
rect 3783 4362 3817 4486
rect 3985 4362 4125 4396
rect 4293 4362 4327 4486
rect 4407 4362 6729 4396
<< viali >>
rect 2995 4362 3029 4396
rect 3669 4362 3703 4396
rect 6729 4362 6763 4396
<< metal1 >>
rect 2816 8648 3597 8682
rect 2530 8577 2590 8590
rect 2530 8525 2534 8577
rect 2586 8568 2590 8577
rect 2586 8534 2668 8568
rect 2816 8547 2850 8648
rect 2986 8534 3038 8540
rect 2586 8525 2590 8534
rect 2530 8512 2590 8525
rect 2543 7822 2577 8512
rect 2887 8494 2986 8522
rect 2986 8476 3038 8482
rect 2507 7788 2577 7822
rect 2534 7631 2586 7637
rect 2507 7588 2534 7622
rect 2534 7573 2586 7579
rect 3563 7448 3597 8648
rect 3818 7631 3870 7637
rect 3818 7573 3870 7579
rect 3827 7526 3861 7573
rect 3815 7480 3873 7526
rect 2507 7388 2577 7422
rect 3563 7407 3817 7448
rect 2543 5561 2577 7388
rect 4091 7230 4239 7260
rect 3783 7025 3817 7165
rect 4091 7148 4125 7230
rect 4081 7142 4133 7148
rect 4081 7084 4133 7090
rect 4237 7025 4295 7189
rect 3783 6984 4295 7025
rect 3815 6822 3873 6984
rect 4075 6790 4081 6804
rect 3871 6760 4081 6790
rect 4075 6752 4081 6760
rect 4133 6752 4139 6804
rect 3783 6412 3817 6512
rect 3871 6490 3905 6502
rect 3783 6378 4019 6412
rect 3653 6306 3659 6315
rect 3460 6272 3659 6306
rect 3653 6263 3659 6272
rect 3711 6263 3717 6315
rect 3494 6164 3873 6210
rect 3563 5832 3817 5867
rect 3865 5832 3951 5874
rect 2534 5555 2586 5561
rect 3460 5506 3500 5552
rect 2534 5497 2586 5503
rect 2893 4510 2933 4538
rect 2893 4476 3225 4510
rect 3563 4471 3597 5832
rect 3660 5555 3712 5561
rect 3815 5546 3873 5552
rect 3712 5512 3873 5546
rect 3815 5506 3873 5512
rect 3660 5497 3712 5503
rect 3917 5474 3951 5832
rect 3865 5432 3951 5474
rect 3985 5432 4019 6378
rect 4091 6321 4125 6752
rect 4082 6315 4134 6321
rect 4082 6257 4134 6263
rect 4091 5821 4125 6257
rect 4287 5862 6696 5890
rect 4091 5765 4295 5821
rect 4237 5464 4295 5765
rect 4339 5432 4373 5862
rect 3985 5395 4239 5432
rect 4287 5404 4373 5432
rect 4159 5132 4239 5161
rect 4159 4774 4193 5132
rect 4293 4812 4327 5156
rect 4159 4745 4239 4774
rect 3378 4437 3597 4471
rect 6707 4405 6785 4409
rect 2983 4396 3041 4402
rect 3663 4396 3715 4402
rect 2983 4362 2995 4396
rect 3029 4362 3669 4396
rect 3703 4362 3715 4396
rect 2983 4356 3041 4362
rect 3663 4356 3715 4362
rect 6707 4353 6720 4405
rect 6772 4353 6785 4405
rect 6707 4349 6785 4353
<< via1 >>
rect 2534 8525 2586 8577
rect 2986 8482 3038 8534
rect 2534 7579 2586 7631
rect 3818 7579 3870 7631
rect 4081 7090 4133 7142
rect 4081 6752 4133 6804
rect 3659 6263 3711 6315
rect 2534 5503 2586 5555
rect 3660 5503 3712 5555
rect 4082 6263 4134 6315
rect 6720 4396 6772 4405
rect 6720 4362 6729 4396
rect 6729 4362 6763 4396
rect 6763 4362 6772 4396
rect 6720 4353 6772 4362
<< metal2 >>
rect 2530 8581 2590 8590
rect 2530 8512 2590 8521
rect 2986 8534 3038 8540
rect 6747 8525 6756 8538
rect 3038 8491 6756 8525
rect 2986 8476 3038 8482
rect 6747 8478 6756 8491
rect 6816 8478 6825 8538
rect 3818 7631 3870 7637
rect 2528 7579 2534 7631
rect 2586 7622 2592 7631
rect 2586 7588 3818 7622
rect 2586 7579 2592 7588
rect 3818 7573 3870 7579
rect 4075 7090 4081 7142
rect 4133 7090 4139 7142
rect 4092 6810 4122 7090
rect 4081 6804 4133 6810
rect 4081 6746 4133 6752
rect 3659 6315 3711 6321
rect 4076 6306 4082 6315
rect 3711 6272 4082 6306
rect 4076 6263 4082 6272
rect 4134 6263 4140 6315
rect 3659 6257 3711 6263
rect 3660 5555 3712 5561
rect 2528 5503 2534 5555
rect 2586 5546 2592 5555
rect 2586 5512 3660 5546
rect 2586 5503 2592 5512
rect 3660 5497 3712 5503
rect 6707 4349 6716 4409
rect 6776 4349 6785 4409
<< via2 >>
rect 2530 8577 2590 8581
rect 2530 8525 2534 8577
rect 2534 8525 2586 8577
rect 2586 8525 2590 8577
rect 2530 8521 2590 8525
rect 6756 8478 6816 8538
rect 6716 4405 6776 4409
rect 6716 4353 6720 4405
rect 6720 4353 6772 4405
rect 6772 4353 6776 4405
rect 6716 4349 6776 4353
<< metal3 >>
rect 2525 8581 2595 8586
rect 2525 8521 2530 8581
rect 2590 8521 2777 8581
rect 2525 8516 2595 8521
rect 2717 8422 2777 8521
rect 6751 8538 6821 8543
rect 6751 8478 6756 8538
rect 6816 8478 7081 8538
rect 6751 8473 6821 8478
rect 6714 4583 6778 4589
rect 6714 4513 6778 4519
rect 6716 4414 6776 4513
rect 6711 4409 6781 4414
rect 6711 4349 6716 4409
rect 6776 4349 6781 4409
rect 6711 4344 6781 4349
<< via3 >>
rect 6714 4519 6778 4583
<< metal4 >>
rect 6416 8025 6851 8106
rect 6713 4583 6779 4584
rect 6713 4581 6714 4583
rect 6420 4521 6714 4581
rect 6713 4519 6714 4521
rect 6778 4519 6779 4583
rect 6713 4518 6779 4519
use sky130_fd_pr__cap_mim_m3_1_BNHTNG  sky130_fd_pr__cap_mim_m3_1_BNHTNG_0
timestamp 1728522838
transform 0 1 4547 1 0 6512
box -2186 -2040 2186 2040
use sky130_fd_pr__nfet_01v8_84Z3BM  sky130_fd_pr__nfet_01v8_84Z3BM_0
timestamp 1728500067
transform 1 0 3844 0 1 7329
box -211 -329 211 329
use sky130_fd_pr__pfet_01v8_ZMS3C4  sky130_fd_pr__pfet_01v8_ZMS3C4_0
timestamp 1728002984
transform 0 1 3349 -1 0 6522
box -2196 -284 2196 284
use sky130_fd_pr__cap_mim_m3_1_EYXEMC  XC2
timestamp 1728608927
transform 0 -1 7215 1 0 7512
box -1186 -540 1186 540
use sky130_fd_pr__nfet_01v8_QXQH2M  XM2
timestamp 1727994832
transform 0 1 2786 -1 0 6522
box -2196 -279 2196 279
use sky130_fd_pr__nfet_01v8_84Z3BM  XM4
timestamp 1728500067
transform 1 0 3844 0 1 6013
box -211 -329 211 329
use sky130_fd_pr__nfet_01v8_BBX9LZ  XM5
timestamp 1727994832
transform 1 0 3844 0 1 5005
box -211 -679 211 679
use sky130_fd_pr__pfet_01v8_LJP3BL  XM6
timestamp 1728501028
transform 1 0 4266 0 1 7344
box -211 -334 211 334
use sky130_fd_pr__nfet_01v8_84Z3BM  XM7
timestamp 1728500067
transform -1 0 3844 0 1 6671
box -211 -329 211 329
use sky130_fd_pr__pfet_01v8_MGSVTG  XM8
timestamp 1728501028
transform 1 0 4266 0 1 6326
box -211 -684 211 684
use sky130_fd_pr__nfet_01v8_84Z3BM  XM9
timestamp 1728500067
transform -1 0 4266 0 1 5313
box -211 -329 211 329
use sky130_fd_pr__nfet_01v8_84Z3BM  XM10
timestamp 1728500067
transform 1 0 4266 0 1 4655
box -211 -329 211 329
<< labels >>
flabel locali s 2543 4326 2613 4326 0 FreeSans 480 0 0 0 GND
port 0 nsew
flabel locali s 3563 8718 3633 8718 0 FreeSans 480 0 0 0 VDD
port 1 nsew
flabel metal1 s 2507 7788 2507 7822 0 FreeSans 480 0 0 0 Iin
port 2 nsew
flabel metal1 s 2507 7588 2507 7622 0 FreeSans 480 0 0 0 Vlky
port 3 nsew
flabel metal1 s 2507 7388 2507 7422 0 FreeSans 480 0 0 0 Vb
port 4 nsew
<< end >>
