magic
tech sky130B
magscale 1 2
timestamp 1728498447
<< nwell >>
rect -696 -269 696 269
<< pmos >>
rect -500 -50 500 50
<< pdiff >>
rect -558 38 -500 50
rect -558 -38 -546 38
rect -512 -38 -500 38
rect -558 -50 -500 -38
rect 500 38 558 50
rect 500 -38 512 38
rect 546 -38 558 38
rect 500 -50 558 -38
<< pdiffc >>
rect -546 -38 -512 38
rect 512 -38 546 38
<< nsubdiff >>
rect -660 199 -564 233
rect 564 199 660 233
rect -660 137 -626 199
rect 626 137 660 199
rect -660 -199 -626 -137
rect 626 -199 660 -137
rect -660 -233 -564 -199
rect 564 -233 660 -199
<< nsubdiffcont >>
rect -564 199 564 233
rect -660 -137 -626 137
rect 626 -137 660 137
rect -564 -233 564 -199
<< poly >>
rect -500 131 500 147
rect -500 97 -484 131
rect 484 97 500 131
rect -500 50 500 97
rect -500 -97 500 -50
rect -500 -131 -484 -97
rect 484 -131 500 -97
rect -500 -147 500 -131
<< polycont >>
rect -484 97 484 131
rect -484 -131 484 -97
<< locali >>
rect -660 199 -564 233
rect 564 199 660 233
rect -660 137 -626 199
rect 626 137 660 199
rect -500 97 -484 131
rect 484 97 500 131
rect -546 38 -512 54
rect -546 -54 -512 -38
rect 512 38 546 54
rect 512 -54 546 -38
rect -500 -131 -484 -97
rect 484 -131 500 -97
rect -660 -199 -626 -137
rect 626 -199 660 -137
rect -660 -233 -564 -199
rect 564 -233 660 -199
<< viali >>
rect -484 97 484 131
rect -546 -38 -512 38
rect 512 -38 546 38
rect -484 -131 484 -97
<< metal1 >>
rect -496 131 496 137
rect -496 97 -484 131
rect 484 97 496 131
rect -496 91 496 97
rect -552 38 -506 50
rect -552 -38 -546 38
rect -512 -38 -506 38
rect -552 -50 -506 -38
rect 506 38 552 50
rect 506 -38 512 38
rect 546 -38 552 38
rect 506 -50 552 -38
rect -496 -97 496 -91
rect -496 -131 -484 -97
rect 484 -131 496 -97
rect -496 -137 496 -131
<< properties >>
string FIXED_BBOX -643 -216 643 216
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.5 l 5.0 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
