magic
tech sky130B
magscale 1 2
timestamp 1727994832
<< metal3 >>
rect -1186 512 1186 540
rect -1186 -512 1102 512
rect 1166 -512 1186 512
rect -1186 -540 1186 -512
<< via3 >>
rect 1102 -512 1166 512
<< mimcap >>
rect -1146 460 854 500
rect -1146 -460 -1106 460
rect 814 -460 854 460
rect -1146 -500 854 -460
<< mimcapcontact >>
rect -1106 -460 814 460
<< metal4 >>
rect 1086 512 1182 528
rect -1107 460 815 461
rect -1107 -460 -1106 460
rect 814 -460 815 460
rect -1107 -461 815 -460
rect 1086 -512 1102 512
rect 1166 -512 1182 512
rect 1086 -528 1182 -512
<< properties >>
string FIXED_BBOX -1186 -540 894 540
string gencell sky130_fd_pr__cap_mim_m3_1
string library sky130
string parameters w 10.0 l 5.0 val 105.7 carea 2.00 cperi 0.19 nx 1 ny 1 dummy 0 square 0 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1 ccov 100
<< end >>
