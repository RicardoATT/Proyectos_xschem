** sch_path: /home/ricardo/RATT_repos/Proyectos_xschem/delay/delay_test.sch
**.subckt delay_test
V1 VDD GND 1.8
x1 VDD vin delay GND delay
V2 vin GND PULSE(0 1.8 1n 1n 1n 5n 15n 200)
**** begin user architecture code

.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ricardo/pdk/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/ricardo/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ricardo/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ricardo/pdk/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice


** opencircuitdesign pdks install
.inc /home/ricardo/pdk/sky130B/libs.tech/ngspice/rram_v0.spice



.param Lp_delay=2.15
.param Wp_delay=0.45
.param Ln_delay=2.15
.param Wn_delay=0.45
.control
  save all
  tran 0.1n 1u
  write delay_test.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  /home/ricardo/RATT_repos/Proyectos_xschem/delay/delay.sym # of pins=4
** sym_path: /home/ricardo/RATT_repos/Proyectos_xschem/delay/delay.sym
** sch_path: /home/ricardo/RATT_repos/Proyectos_xschem/delay/delay.sch
.subckt delay VDD Vin Vout GND
*.ipin Vin
*.opin Vout
*.iopin VDD
*.iopin GND
XM1 net1 Vin VDD VDD sky130_fd_pr__pfet_01v8 L={Lp_delay} W={Wp_delay} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 Vin GND GND sky130_fd_pr__nfet_01v8 L={Ln_delay} W={Wn_delay} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 net1 VDD VDD sky130_fd_pr__pfet_01v8 L={Lp_delay} W={Wp_delay} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L={Ln_delay} W={Wn_delay} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM5 net3 net2 VDD VDD sky130_fd_pr__pfet_01v8 L={Lp_delay} W={Wp_delay} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM6 net3 net2 GND GND sky130_fd_pr__nfet_01v8 L={Ln_delay} W={Wn_delay} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout net3 VDD VDD sky130_fd_pr__pfet_01v8 L={Lp_delay} W={Wp_delay} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM8 Vout net3 GND GND sky130_fd_pr__nfet_01v8 L={Ln_delay} W={Wn_delay} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
