magic
tech sky130B
magscale 1 2
timestamp 1728522838
<< pwell >>
rect -246 -710 246 710
<< nmos >>
rect -50 -500 50 500
<< ndiff >>
rect -108 488 -50 500
rect -108 -488 -96 488
rect -62 -488 -50 488
rect -108 -500 -50 -488
rect 50 488 108 500
rect 50 -488 62 488
rect 96 -488 108 488
rect 50 -500 108 -488
<< ndiffc >>
rect -96 -488 -62 488
rect 62 -488 96 488
<< psubdiff >>
rect -210 640 -114 674
rect 114 640 210 674
rect -210 578 -176 640
rect 176 578 210 640
rect -210 -640 -176 -578
rect 176 -640 210 -578
rect -210 -674 -114 -640
rect 114 -674 210 -640
<< psubdiffcont >>
rect -114 640 114 674
rect -210 -578 -176 578
rect 176 -578 210 578
rect -114 -674 114 -640
<< poly >>
rect -50 572 50 588
rect -50 538 -34 572
rect 34 538 50 572
rect -50 500 50 538
rect -50 -538 50 -500
rect -50 -572 -34 -538
rect 34 -572 50 -538
rect -50 -588 50 -572
<< polycont >>
rect -34 538 34 572
rect -34 -572 34 -538
<< locali >>
rect -210 640 -114 674
rect 114 640 210 674
rect -210 578 -176 640
rect 176 578 210 640
rect -50 538 -34 572
rect 34 538 50 572
rect -96 488 -62 504
rect -96 -504 -62 -488
rect 62 488 96 504
rect 62 -504 96 -488
rect -50 -572 -34 -538
rect 34 -572 50 -538
rect -210 -640 -176 -578
rect 176 -640 210 -578
rect -210 -674 -114 -640
rect 114 -674 210 -640
<< viali >>
rect -34 538 34 572
rect -96 -488 -62 488
rect 62 -488 96 488
rect -34 -572 34 -538
<< metal1 >>
rect -46 572 46 578
rect -46 538 -34 572
rect 34 538 46 572
rect -46 532 46 538
rect -102 488 -56 500
rect -102 -488 -96 488
rect -62 -488 -56 488
rect -102 -500 -56 -488
rect 56 488 102 500
rect 56 -488 62 488
rect 96 -488 102 488
rect 56 -500 102 -488
rect -46 -538 46 -532
rect -46 -572 -34 -538
rect 34 -572 46 -538
rect -46 -578 46 -572
<< labels >>
flabel metal1 s -82 31 -82 31 0 FreeSans 480 0 0 0 D
port 24 nsew
flabel metal1 s 82 27 82 27 0 FreeSans 480 0 0 0 S
port 25 nsew
flabel metal1 s -1 -554 -1 -554 0 FreeSans 480 0 0 0 G
port 26 nsew
flabel locali s 1 -660 1 -660 0 FreeSans 480 0 0 0 B
port 27 nsew
<< properties >>
string FIXED_BBOX -193 -657 193 657
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 5.0 l 0.5 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
