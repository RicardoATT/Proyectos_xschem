magic
tech sky130B
magscale 1 2
timestamp 1728432946
<< error_s >>
rect 1352 1487 1387 1496
rect 1459 1487 1809 1496
rect 1370 1381 1792 1451
rect 1370 963 1809 1381
rect 1370 893 1792 963
rect 1406 876 1792 893
rect 1423 840 1792 876
<< locali >>
rect 1387 1949 1459 2019
rect 1071 1841 1151 1875
rect 1071 1211 1151 1245
rect 1387 930 1459 963
rect 1387 929 1493 930
rect 1459 823 1493 929
rect 1493 653 1573 687
rect 1387 335 1459 405
<< metal1 >>
rect 1239 1671 1319 1699
rect 1195 1521 1229 1624
rect 1285 1536 1319 1671
rect 1527 1671 1573 1699
rect 1695 1671 1741 1699
rect 1001 1487 1229 1521
rect 1028 1424 1080 1430
rect 1001 1381 1028 1415
rect 1028 1366 1080 1372
rect 1195 1313 1229 1487
rect 1276 1530 1328 1536
rect 1276 1472 1328 1478
rect 1037 1279 1229 1313
rect 1037 963 1071 1279
rect 1285 1241 1319 1472
rect 1527 1430 1561 1671
rect 1617 1536 1651 1624
rect 1608 1530 1660 1536
rect 1608 1472 1660 1478
rect 1707 1521 1741 1671
rect 1707 1487 1845 1521
rect 1518 1424 1570 1430
rect 1518 1366 1570 1372
rect 1527 1303 1561 1366
rect 1707 1303 1741 1487
rect 1527 1275 1573 1303
rect 1239 1213 1319 1241
rect 1695 1103 1741 1303
rect 1617 963 1651 1065
rect 1037 929 1651 963
rect 1001 823 1651 857
rect 1617 721 1651 823
rect 1707 683 1741 1103
rect 1695 655 1741 683
<< via1 >>
rect 1028 1372 1080 1424
rect 1276 1478 1328 1530
rect 1608 1478 1660 1530
rect 1518 1372 1570 1424
<< metal2 >>
rect 1270 1478 1276 1530
rect 1328 1521 1334 1530
rect 1602 1521 1608 1530
rect 1328 1487 1608 1521
rect 1328 1478 1334 1487
rect 1602 1478 1608 1487
rect 1660 1478 1666 1530
rect 1022 1372 1028 1424
rect 1080 1415 1086 1424
rect 1512 1415 1518 1424
rect 1080 1381 1518 1415
rect 1080 1372 1086 1381
rect 1512 1372 1518 1381
rect 1570 1372 1576 1424
use sky130_fd_pr__pfet_01v8_LGS3BL  sky130_fd_pr__pfet_01v8_LGS3BL_0
timestamp 1728430153
transform 1 0 1634 0 1 1735
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_LGS3BL  XM1
timestamp 1728430153
transform 1 0 1212 0 1 1735
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1728430153
transform 1 0 1212 0 1 1172
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 0
transform 1 0 1581 0 1 1159
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_64QSBY  XM4
timestamp 1728430229
transform 1 0 1634 0 1 1172
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_64Z3AY  XM5
timestamp 1728430153
transform 1 0 1634 0 1 614
box -211 -279 211 279
<< labels >>
flabel locali s 1387 335 1459 335 0 FreeSans 480 0 0 0 GND
port 12 nsew
flabel locali s 1387 2019 1459 2019 0 FreeSans 480 0 0 0 VDD
port 13 nsew
flabel metal1 s 1845 1487 1845 1521 0 FreeSans 480 0 0 0 Vout
port 14 nsew
flabel metal1 s 1001 1487 1001 1521 0 FreeSans 480 0 0 0 Ctrl
port 15 nsew
flabel metal1 s 1001 1381 1001 1415 0 FreeSans 480 0 0 0 Vin
port 16 nsew
flabel metal1 s 1001 823 1001 857 0 FreeSans 480 0 0 0 Vbias
port 17 nsew
<< end >>
