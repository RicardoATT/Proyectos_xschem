magic
tech sky130B
magscale 1 2
timestamp 1728085572
<< locali >>
rect 3101 8534 3297 8568
rect 3597 7682 4125 7692
rect 3563 7658 4125 7682
rect 4091 7608 4125 7658
rect 4293 7503 4327 7642
rect 3669 6930 3703 7070
rect 3871 7036 3905 7160
rect 4091 6940 4125 7080
rect 4205 6825 4239 6974
rect 3669 6272 3703 6412
rect 3669 5614 3703 5754
rect 4091 4914 4125 5054
rect 2651 4362 2687 4510
rect 3783 4362 3817 4486
rect 3985 4362 4125 4396
rect 4293 4362 4327 4486
<< viali >>
rect 2995 4362 3029 4396
rect 3669 4362 3703 4396
<< metal1 >>
rect 2816 8648 3597 8682
rect 2816 8547 2850 8648
rect 3563 7448 3597 8648
rect 3815 7480 3873 7571
rect 3563 7407 3817 7448
rect 4091 7230 4239 7260
rect 3783 7025 3817 7165
rect 4091 7148 4125 7230
rect 4081 7142 4133 7148
rect 4081 7084 4133 7090
rect 4237 7025 4295 7189
rect 3783 6984 4295 7025
rect 3815 6822 3873 6984
rect 4075 6790 4081 6804
rect 3871 6760 4081 6790
rect 4075 6752 4081 6760
rect 4133 6752 4139 6804
rect 3783 6412 3817 6512
rect 3871 6490 3905 6502
rect 3783 6378 4019 6412
rect 3653 6306 3659 6315
rect 3460 6272 3659 6306
rect 3653 6263 3659 6272
rect 3711 6263 3717 6315
rect 3494 6164 3873 6210
rect 3563 5832 3817 5867
rect 3865 5832 3951 5874
rect 3460 5506 3500 5552
rect 3563 4471 3597 5832
rect 3815 5506 3873 5597
rect 3917 5474 3951 5832
rect 3865 5432 3951 5474
rect 3985 5432 4019 6378
rect 4091 6321 4125 6752
rect 4082 6315 4134 6321
rect 4082 6257 4134 6263
rect 4091 5821 4125 6257
rect 4287 5862 4373 5890
rect 4091 5765 4295 5821
rect 4237 5464 4295 5765
rect 4339 5432 4373 5862
rect 3985 5395 4239 5432
rect 4287 5404 4373 5432
rect 4159 5132 4239 5161
rect 4159 4774 4193 5132
rect 4293 4812 4327 5156
rect 4159 4745 4239 4774
rect 3378 4437 3597 4471
rect 2983 4396 3041 4402
rect 3663 4396 3715 4402
rect 2983 4362 2995 4396
rect 3029 4362 3669 4396
rect 3703 4362 3715 4396
rect 2983 4356 3041 4362
rect 3663 4356 3715 4362
<< via1 >>
rect 4081 7090 4133 7142
rect 4081 6752 4133 6804
rect 3659 6263 3711 6315
rect 4082 6263 4134 6315
<< metal2 >>
rect 4075 7090 4081 7142
rect 4133 7090 4139 7142
rect 4092 6810 4122 7090
rect 4081 6804 4133 6810
rect 4081 6746 4133 6752
rect 3659 6315 3711 6321
rect 4076 6306 4082 6315
rect 3711 6272 4082 6306
rect 4076 6263 4082 6272
rect 4134 6263 4140 6315
rect 3659 6257 3711 6263
use sky130_fd_pr__cap_mim_m3_1_BNHTNG  sky130_fd_pr__cap_mim_m3_1_BNHTNG_1
timestamp 1728085572
transform 0 -1 13322 1 0 6071
box -2186 -2040 2186 2040
use sky130_fd_pr__nfet_01v8_84Z3BM  sky130_fd_pr__nfet_01v8_84Z3BM_0
timestamp 1727994832
transform 1 0 3844 0 1 7329
box -211 -329 211 329
use sky130_fd_pr__pfet_01v8_ZMS3C4  sky130_fd_pr__pfet_01v8_ZMS3C4_0
timestamp 1728002984
transform 0 1 3349 -1 0 6522
box -2196 -284 2196 284
use sky130_fd_pr__cap_mim_m3_1_EYXEMC  XC2
timestamp 1727994832
transform 0 -1 7215 1 0 7512
box -1186 -540 1186 540
use sky130_fd_pr__nfet_01v8_QXQH2M  XM2
timestamp 1727994832
transform 0 1 2786 -1 0 6522
box -2196 -279 2196 279
use sky130_fd_pr__nfet_01v8_84Z3BM  XM4
timestamp 1727994832
transform 1 0 3844 0 1 6013
box -211 -329 211 329
use sky130_fd_pr__nfet_01v8_BBX9LZ  XM5
timestamp 1727994832
transform 1 0 3844 0 1 5005
box -211 -679 211 679
use sky130_fd_pr__pfet_01v8_LJP3BL  XM6
timestamp 1727994832
transform 1 0 4266 0 1 7344
box -211 -334 211 334
use sky130_fd_pr__nfet_01v8_84Z3BM  XM7
timestamp 1727994832
transform -1 0 3844 0 1 6671
box -211 -329 211 329
use sky130_fd_pr__pfet_01v8_MGSVTG  XM8
timestamp 1727994832
transform 1 0 4266 0 1 6326
box -211 -684 211 684
use sky130_fd_pr__nfet_01v8_84Z3BM  XM9
timestamp 1727994832
transform -1 0 4266 0 1 5313
box -211 -329 211 329
use sky130_fd_pr__nfet_01v8_84Z3BM  XM10
timestamp 1727994832
transform 1 0 4266 0 1 4655
box -211 -329 211 329
<< end >>
