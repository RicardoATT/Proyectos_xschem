magic
tech sky130B
magscale 1 2
timestamp 1729119800
<< error_p >>
rect -605 172 -547 178
rect -413 172 -355 178
rect -221 172 -163 178
rect -29 172 29 178
rect 163 172 221 178
rect 355 172 413 178
rect 547 172 605 178
rect -605 138 -593 172
rect -413 138 -401 172
rect -221 138 -209 172
rect -29 138 -17 172
rect 163 138 175 172
rect 355 138 367 172
rect 547 138 559 172
rect -605 132 -547 138
rect -413 132 -355 138
rect -221 132 -163 138
rect -29 132 29 138
rect 163 132 221 138
rect 355 132 413 138
rect 547 132 605 138
rect -701 -138 -643 -132
rect -509 -138 -451 -132
rect -317 -138 -259 -132
rect -125 -138 -67 -132
rect 67 -138 125 -132
rect 259 -138 317 -132
rect 451 -138 509 -132
rect 643 -138 701 -132
rect -701 -172 -689 -138
rect -509 -172 -497 -138
rect -317 -172 -305 -138
rect -125 -172 -113 -138
rect 67 -172 79 -138
rect 259 -172 271 -138
rect 451 -172 463 -138
rect 643 -172 655 -138
rect -701 -178 -643 -172
rect -509 -178 -451 -172
rect -317 -178 -259 -172
rect -125 -178 -67 -172
rect 67 -178 125 -172
rect 259 -178 317 -172
rect 451 -178 509 -172
rect 643 -178 701 -172
<< pwell >>
rect -887 -310 887 310
<< nmos >>
rect -687 -100 -657 100
rect -591 -100 -561 100
rect -495 -100 -465 100
rect -399 -100 -369 100
rect -303 -100 -273 100
rect -207 -100 -177 100
rect -111 -100 -81 100
rect -15 -100 15 100
rect 81 -100 111 100
rect 177 -100 207 100
rect 273 -100 303 100
rect 369 -100 399 100
rect 465 -100 495 100
rect 561 -100 591 100
rect 657 -100 687 100
<< ndiff >>
rect -749 88 -687 100
rect -749 -88 -737 88
rect -703 -88 -687 88
rect -749 -100 -687 -88
rect -657 88 -591 100
rect -657 -88 -641 88
rect -607 -88 -591 88
rect -657 -100 -591 -88
rect -561 88 -495 100
rect -561 -88 -545 88
rect -511 -88 -495 88
rect -561 -100 -495 -88
rect -465 88 -399 100
rect -465 -88 -449 88
rect -415 -88 -399 88
rect -465 -100 -399 -88
rect -369 88 -303 100
rect -369 -88 -353 88
rect -319 -88 -303 88
rect -369 -100 -303 -88
rect -273 88 -207 100
rect -273 -88 -257 88
rect -223 -88 -207 88
rect -273 -100 -207 -88
rect -177 88 -111 100
rect -177 -88 -161 88
rect -127 -88 -111 88
rect -177 -100 -111 -88
rect -81 88 -15 100
rect -81 -88 -65 88
rect -31 -88 -15 88
rect -81 -100 -15 -88
rect 15 88 81 100
rect 15 -88 31 88
rect 65 -88 81 88
rect 15 -100 81 -88
rect 111 88 177 100
rect 111 -88 127 88
rect 161 -88 177 88
rect 111 -100 177 -88
rect 207 88 273 100
rect 207 -88 223 88
rect 257 -88 273 88
rect 207 -100 273 -88
rect 303 88 369 100
rect 303 -88 319 88
rect 353 -88 369 88
rect 303 -100 369 -88
rect 399 88 465 100
rect 399 -88 415 88
rect 449 -88 465 88
rect 399 -100 465 -88
rect 495 88 561 100
rect 495 -88 511 88
rect 545 -88 561 88
rect 495 -100 561 -88
rect 591 88 657 100
rect 591 -88 607 88
rect 641 -88 657 88
rect 591 -100 657 -88
rect 687 88 749 100
rect 687 -88 703 88
rect 737 -88 749 88
rect 687 -100 749 -88
<< ndiffc >>
rect -737 -88 -703 88
rect -641 -88 -607 88
rect -545 -88 -511 88
rect -449 -88 -415 88
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect 415 -88 449 88
rect 511 -88 545 88
rect 607 -88 641 88
rect 703 -88 737 88
<< psubdiff >>
rect -851 240 -755 274
rect 755 240 851 274
rect -851 178 -817 240
rect 817 178 851 240
rect -851 -240 -817 -178
rect 817 -240 851 -178
rect -851 -274 -755 -240
rect 755 -274 851 -240
<< psubdiffcont >>
rect -755 240 755 274
rect -851 -178 -817 178
rect 817 -178 851 178
rect -755 -274 755 -240
<< poly >>
rect -609 172 -543 188
rect -609 138 -593 172
rect -559 138 -543 172
rect -687 100 -657 126
rect -609 122 -543 138
rect -417 172 -351 188
rect -417 138 -401 172
rect -367 138 -351 172
rect -591 100 -561 122
rect -495 100 -465 126
rect -417 122 -351 138
rect -225 172 -159 188
rect -225 138 -209 172
rect -175 138 -159 172
rect -399 100 -369 122
rect -303 100 -273 126
rect -225 122 -159 138
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -207 100 -177 122
rect -111 100 -81 126
rect -33 122 33 138
rect 159 172 225 188
rect 159 138 175 172
rect 209 138 225 172
rect -15 100 15 122
rect 81 100 111 126
rect 159 122 225 138
rect 351 172 417 188
rect 351 138 367 172
rect 401 138 417 172
rect 177 100 207 122
rect 273 100 303 126
rect 351 122 417 138
rect 543 172 609 188
rect 543 138 559 172
rect 593 138 609 172
rect 369 100 399 122
rect 465 100 495 126
rect 543 122 609 138
rect 561 100 591 122
rect 657 100 687 126
rect -687 -122 -657 -100
rect -705 -138 -639 -122
rect -591 -126 -561 -100
rect -495 -122 -465 -100
rect -705 -172 -689 -138
rect -655 -172 -639 -138
rect -705 -188 -639 -172
rect -513 -138 -447 -122
rect -399 -126 -369 -100
rect -303 -122 -273 -100
rect -513 -172 -497 -138
rect -463 -172 -447 -138
rect -513 -188 -447 -172
rect -321 -138 -255 -122
rect -207 -126 -177 -100
rect -111 -122 -81 -100
rect -321 -172 -305 -138
rect -271 -172 -255 -138
rect -321 -188 -255 -172
rect -129 -138 -63 -122
rect -15 -126 15 -100
rect 81 -122 111 -100
rect -129 -172 -113 -138
rect -79 -172 -63 -138
rect -129 -188 -63 -172
rect 63 -138 129 -122
rect 177 -126 207 -100
rect 273 -122 303 -100
rect 63 -172 79 -138
rect 113 -172 129 -138
rect 63 -188 129 -172
rect 255 -138 321 -122
rect 369 -126 399 -100
rect 465 -122 495 -100
rect 255 -172 271 -138
rect 305 -172 321 -138
rect 255 -188 321 -172
rect 447 -138 513 -122
rect 561 -126 591 -100
rect 657 -122 687 -100
rect 447 -172 463 -138
rect 497 -172 513 -138
rect 447 -188 513 -172
rect 639 -138 705 -122
rect 639 -172 655 -138
rect 689 -172 705 -138
rect 639 -188 705 -172
<< polycont >>
rect -593 138 -559 172
rect -401 138 -367 172
rect -209 138 -175 172
rect -17 138 17 172
rect 175 138 209 172
rect 367 138 401 172
rect 559 138 593 172
rect -689 -172 -655 -138
rect -497 -172 -463 -138
rect -305 -172 -271 -138
rect -113 -172 -79 -138
rect 79 -172 113 -138
rect 271 -172 305 -138
rect 463 -172 497 -138
rect 655 -172 689 -138
<< locali >>
rect -851 240 -755 274
rect 755 240 851 274
rect -851 178 -817 240
rect 817 178 851 240
rect -609 138 -593 172
rect -559 138 -543 172
rect -417 138 -401 172
rect -367 138 -351 172
rect -225 138 -209 172
rect -175 138 -159 172
rect -33 138 -17 172
rect 17 138 33 172
rect 159 138 175 172
rect 209 138 225 172
rect 351 138 367 172
rect 401 138 417 172
rect 543 138 559 172
rect 593 138 609 172
rect -737 88 -703 104
rect -737 -104 -703 -88
rect -641 88 -607 104
rect -641 -104 -607 -88
rect -545 88 -511 104
rect -545 -104 -511 -88
rect -449 88 -415 104
rect -449 -104 -415 -88
rect -353 88 -319 104
rect -353 -104 -319 -88
rect -257 88 -223 104
rect -257 -104 -223 -88
rect -161 88 -127 104
rect -161 -104 -127 -88
rect -65 88 -31 104
rect -65 -104 -31 -88
rect 31 88 65 104
rect 31 -104 65 -88
rect 127 88 161 104
rect 127 -104 161 -88
rect 223 88 257 104
rect 223 -104 257 -88
rect 319 88 353 104
rect 319 -104 353 -88
rect 415 88 449 104
rect 415 -104 449 -88
rect 511 88 545 104
rect 511 -104 545 -88
rect 607 88 641 104
rect 607 -104 641 -88
rect 703 88 737 104
rect 703 -104 737 -88
rect -705 -172 -689 -138
rect -655 -172 -639 -138
rect -513 -172 -497 -138
rect -463 -172 -447 -138
rect -321 -172 -305 -138
rect -271 -172 -255 -138
rect -129 -172 -113 -138
rect -79 -172 -63 -138
rect 63 -172 79 -138
rect 113 -172 129 -138
rect 255 -172 271 -138
rect 305 -172 321 -138
rect 447 -172 463 -138
rect 497 -172 513 -138
rect 639 -172 655 -138
rect 689 -172 705 -138
rect -851 -240 -817 -178
rect 817 -240 851 -178
rect -851 -274 -755 -240
rect 755 -274 851 -240
<< viali >>
rect -593 138 -559 172
rect -401 138 -367 172
rect -209 138 -175 172
rect -17 138 17 172
rect 175 138 209 172
rect 367 138 401 172
rect 559 138 593 172
rect -737 -88 -703 88
rect -641 -88 -607 88
rect -545 -88 -511 88
rect -449 -88 -415 88
rect -353 -88 -319 88
rect -257 -88 -223 88
rect -161 -88 -127 88
rect -65 -88 -31 88
rect 31 -88 65 88
rect 127 -88 161 88
rect 223 -88 257 88
rect 319 -88 353 88
rect 415 -88 449 88
rect 511 -88 545 88
rect 607 -88 641 88
rect 703 -88 737 88
rect -689 -172 -655 -138
rect -497 -172 -463 -138
rect -305 -172 -271 -138
rect -113 -172 -79 -138
rect 79 -172 113 -138
rect 271 -172 305 -138
rect 463 -172 497 -138
rect 655 -172 689 -138
<< metal1 >>
rect -605 172 -547 178
rect -605 138 -593 172
rect -559 138 -547 172
rect -605 132 -547 138
rect -413 172 -355 178
rect -413 138 -401 172
rect -367 138 -355 172
rect -413 132 -355 138
rect -221 172 -163 178
rect -221 138 -209 172
rect -175 138 -163 172
rect -221 132 -163 138
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect 163 172 221 178
rect 163 138 175 172
rect 209 138 221 172
rect 163 132 221 138
rect 355 172 413 178
rect 355 138 367 172
rect 401 138 413 172
rect 355 132 413 138
rect 547 172 605 178
rect 547 138 559 172
rect 593 138 605 172
rect 547 132 605 138
rect -743 88 -697 100
rect -743 -88 -737 88
rect -703 -88 -697 88
rect -743 -100 -697 -88
rect -647 88 -601 100
rect -647 -88 -641 88
rect -607 -88 -601 88
rect -647 -100 -601 -88
rect -551 88 -505 100
rect -551 -88 -545 88
rect -511 -88 -505 88
rect -551 -100 -505 -88
rect -455 88 -409 100
rect -455 -88 -449 88
rect -415 -88 -409 88
rect -455 -100 -409 -88
rect -359 88 -313 100
rect -359 -88 -353 88
rect -319 -88 -313 88
rect -359 -100 -313 -88
rect -263 88 -217 100
rect -263 -88 -257 88
rect -223 -88 -217 88
rect -263 -100 -217 -88
rect -167 88 -121 100
rect -167 -88 -161 88
rect -127 -88 -121 88
rect -167 -100 -121 -88
rect -71 88 -25 100
rect -71 -88 -65 88
rect -31 -88 -25 88
rect -71 -100 -25 -88
rect 25 88 71 100
rect 25 -88 31 88
rect 65 -88 71 88
rect 25 -100 71 -88
rect 121 88 167 100
rect 121 -88 127 88
rect 161 -88 167 88
rect 121 -100 167 -88
rect 217 88 263 100
rect 217 -88 223 88
rect 257 -88 263 88
rect 217 -100 263 -88
rect 313 88 359 100
rect 313 -88 319 88
rect 353 -88 359 88
rect 313 -100 359 -88
rect 409 88 455 100
rect 409 -88 415 88
rect 449 -88 455 88
rect 409 -100 455 -88
rect 505 88 551 100
rect 505 -88 511 88
rect 545 -88 551 88
rect 505 -100 551 -88
rect 601 88 647 100
rect 601 -88 607 88
rect 641 -88 647 88
rect 601 -100 647 -88
rect 697 88 743 100
rect 697 -88 703 88
rect 737 -88 743 88
rect 697 -100 743 -88
rect -701 -138 -643 -132
rect -701 -172 -689 -138
rect -655 -172 -643 -138
rect -701 -178 -643 -172
rect -509 -138 -451 -132
rect -509 -172 -497 -138
rect -463 -172 -451 -138
rect -509 -178 -451 -172
rect -317 -138 -259 -132
rect -317 -172 -305 -138
rect -271 -172 -259 -138
rect -317 -178 -259 -172
rect -125 -138 -67 -132
rect -125 -172 -113 -138
rect -79 -172 -67 -138
rect -125 -178 -67 -172
rect 67 -138 125 -132
rect 67 -172 79 -138
rect 113 -172 125 -138
rect 67 -178 125 -172
rect 259 -138 317 -132
rect 259 -172 271 -138
rect 305 -172 317 -138
rect 259 -178 317 -172
rect 451 -138 509 -132
rect 451 -172 463 -138
rect 497 -172 509 -138
rect 451 -178 509 -172
rect 643 -138 701 -132
rect 643 -172 655 -138
rect 689 -172 701 -138
rect 643 -178 701 -172
<< labels >>
flabel metal1 s -576 155 -576 155 0 FreeSans 480 0 0 0 G
port 0 nsew
flabel metal1 s -720 0 -720 0 0 FreeSans 480 0 0 0 D
port 1 nsew
flabel metal1 s -624 -2 -624 -2 0 FreeSans 480 0 0 0 S
port 2 nsew
flabel locali s -11 -257 -11 -257 0 FreeSans 480 0 0 0 B
port 3 nsew
<< properties >>
string FIXED_BBOX -834 -257 834 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 15 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
