magic
tech sky130B
magscale 1 2
timestamp 1728442182
<< locali >>
rect -4842 4458 -4808 4551
rect -5172 4378 -5092 4412
rect -5546 4238 -5439 4240
rect -5634 4134 -5600 4226
rect -5546 4206 -5434 4238
rect -5634 4100 -5494 4134
rect -5468 4108 -5434 4206
rect -4590 4090 -4556 4230
rect -5916 3992 -5836 4026
rect -4704 3911 -4590 3945
rect -5209 1652 -4872 1686
<< metal1 >>
rect -5882 4548 -4922 4582
rect -5882 4408 -5848 4548
rect -5774 4446 -5234 4480
rect -5882 4379 -5836 4408
rect -5654 4380 -5648 4408
rect -5959 4249 -5907 4255
rect -5959 4191 -5907 4197
rect -5950 1661 -5916 4191
rect -5688 4022 -5654 4330
rect -5574 4255 -5540 4446
rect -5360 4380 -5354 4408
rect -5414 4340 -5360 4346
rect -5414 4318 -5354 4340
rect -5583 4249 -5531 4255
rect -5583 4191 -5531 4197
rect -5714 3994 -5654 4022
rect -5414 4004 -5380 4318
rect -4956 4230 -4922 4548
rect -4670 4392 -4556 4458
rect -4780 4230 -4732 4333
rect -4956 4196 -4732 4230
rect -4780 4028 -4732 4196
rect -4815 4022 -4732 4028
rect -5326 3991 -4814 4022
rect -4805 3991 -4732 4022
rect -5326 3988 -4732 3991
rect -4828 3982 -4766 3988
rect -4886 3932 -4873 3941
rect -4905 3926 -4853 3932
rect -4800 3924 -4766 3982
rect -4713 3926 -4661 3932
rect -4905 3868 -4853 3874
rect -4713 3868 -4661 3874
rect -4992 1900 -4958 1953
rect -4800 1900 -4766 1953
rect -4992 1894 -4930 1900
rect -4800 1894 -4763 1900
rect -4992 1860 -4718 1894
rect -5986 1627 -5916 1661
rect -5959 1593 -5907 1599
rect -5986 1550 -5959 1584
rect -4921 1541 -4915 1593
rect -4863 1584 -4857 1593
rect -4863 1550 -4714 1584
rect -4863 1541 -4857 1550
rect -5959 1535 -5907 1541
rect -5986 1473 -5916 1507
rect -5950 990 -5916 1473
rect -5429 1458 -5423 1510
rect -5371 1458 -5365 1510
rect -5073 1417 -5009 1522
rect -4590 1512 -4556 4392
rect -4670 1484 -4556 1512
rect -5762 1365 -5756 1417
rect -5704 1365 -5698 1417
rect -5073 1365 -5064 1417
rect -5012 1365 -5009 1417
rect -5073 1359 -5009 1365
rect -4792 1134 -4758 1227
rect -4792 1100 -4520 1134
rect -5950 984 -5752 990
rect -5950 950 -5336 984
rect -5950 944 -5752 950
<< via1 >>
rect -5959 4197 -5907 4249
rect -5583 4197 -5531 4249
rect -4905 3874 -4853 3926
rect -4713 3874 -4661 3926
rect -5959 1541 -5907 1593
rect -4915 1541 -4863 1593
rect -5423 1458 -5371 1510
rect -5756 1365 -5704 1417
rect -5064 1365 -5012 1417
<< metal2 >>
rect -5965 4197 -5959 4249
rect -5907 4240 -5901 4249
rect -5589 4240 -5583 4249
rect -5907 4206 -5583 4240
rect -5907 4197 -5901 4206
rect -5589 4197 -5583 4206
rect -5531 4197 -5525 4249
rect -4911 3874 -4905 3926
rect -4853 3914 -4847 3926
rect -4719 3914 -4713 3926
rect -4853 3886 -4713 3914
rect -4853 3874 -4847 3886
rect -4719 3874 -4713 3886
rect -4661 3874 -4655 3926
rect -4915 1593 -4863 1599
rect -5965 1541 -5959 1593
rect -5907 1584 -5901 1593
rect -5907 1550 -4915 1584
rect -5907 1541 -5901 1550
rect -4915 1535 -4863 1541
rect -5423 1510 -5371 1516
rect -5079 1507 -5002 1516
rect -5371 1461 -5002 1507
rect -5423 1452 -5371 1458
rect -5079 1449 -5002 1461
rect -5756 1417 -5704 1423
rect -5070 1414 -5064 1417
rect -5704 1368 -5064 1414
rect -5070 1365 -5064 1368
rect -5012 1365 -5006 1417
rect -5756 1359 -5704 1365
use sky130_fd_pr__nfet_01v8_P46M8Q  sky130_fd_pr__nfet_01v8_P46M8Q_0
timestamp 1728435493
transform 1 0 -5263 0 1 4394
box -241 -224 241 224
use sky130_fd_pr__nfet_01v8_X2WNKZ  sky130_fd_pr__nfet_01v8_X2WNKZ_0
timestamp 1728435493
transform -1 0 -5353 0 1 2491
box -211 -1679 211 1679
use sky130_fd_pr_reram__reram_cell  sky130_fd_pr_reram__reram_cell_0
timestamp 1727988820
transform 1 0 -5041 0 1 1484
box -38 -38 38 38
use sky130_fd_pr__nfet_01v8_P46M8Q  XM1
timestamp 1728435493
transform 1 0 -5745 0 1 4394
box -241 -224 241 224
use sky130_fd_pr__nfet_01v8_X2WNKZ  XM2
timestamp 1728435493
transform -1 0 -5775 0 1 2491
box -211 -1679 211 1679
use sky130_fd_pr__pfet_01v8_UGKMGH  XM5
timestamp 1728435493
transform 1 0 -4831 0 1 2941
box -311 -1219 311 1219
use sky130_fd_pr__pfet_01v8_UAJFQ5  XM6
timestamp 1728435493
transform -1 0 -4756 0 1 4389
box -236 -229 236 229
use sky130_fd_pr__nfet_01v8_84QSGM  XM7
timestamp 1728435493
transform -1 0 -4731 0 -1 1393
box -211 -329 211 329
<< end >>
