magic
tech sky130B
magscale 1 2
timestamp 1728343558
<< locali >>
rect 236 1372 308 1408
rect 202 1338 342 1372
rect -114 1230 34 1264
rect -114 710 34 744
rect 202 538 342 572
rect 308 432 342 538
rect 308 262 448 296
rect 236 54 308 124
<< metal1 >>
rect 88 1170 168 1198
rect 32 812 90 1129
rect -150 778 90 812
rect -114 572 -80 778
rect 32 772 90 778
rect 134 1020 168 1170
rect 376 1170 422 1198
rect 544 1170 590 1198
rect 245 1029 297 1035
rect 134 986 245 1020
rect 134 740 168 986
rect 245 971 297 977
rect 244 923 296 929
rect 244 865 296 871
rect 88 712 168 740
rect 253 572 287 865
rect -114 538 287 572
rect 376 740 410 1170
rect 466 1035 500 1123
rect 457 1029 509 1035
rect 457 971 509 977
rect 457 923 509 929
rect 457 865 509 871
rect 466 778 500 865
rect 556 740 590 1170
rect 376 646 422 740
rect 544 712 590 740
rect 544 678 694 712
rect 544 650 590 678
rect 376 500 410 646
rect -150 466 410 500
rect -150 324 512 370
rect 556 292 590 650
rect 544 262 590 292
<< via1 >>
rect 245 977 297 1029
rect 244 871 296 923
rect 457 977 509 1029
rect 457 871 509 923
<< metal2 >>
rect 239 977 245 1029
rect 297 1020 303 1029
rect 451 1020 457 1029
rect 297 986 457 1020
rect 297 977 303 986
rect 451 977 457 986
rect 509 977 515 1029
rect 238 871 244 923
rect 296 914 302 923
rect 451 914 457 923
rect 296 880 457 914
rect 296 871 302 880
rect 451 871 457 880
rect 509 871 515 923
use sky130_fd_pr__nfet_01v8_DR7ETE  sky130_fd_pr__nfet_01v8_DR7ETE_0
timestamp 1728341492
transform 1 0 61 0 1 726
box -211 -224 211 224
use sky130_fd_pr__pfet_01v8_2779BZ  sky130_fd_pr__pfet_01v8_2779BZ_0
timestamp 1728341492
transform 1 0 61 0 1 1179
box -211 -229 211 229
use sky130_fd_pr__pfet_01v8_2779BZ  XM3
timestamp 1728341492
transform 1 0 483 0 1 1179
box -211 -229 211 229
use sky130_fd_pr__nfet_01v8_DR7ETE  XM4
timestamp 1728341492
transform -1 0 483 0 1 726
box -211 -224 211 224
use sky130_fd_pr__nfet_01v8_DR7ETE  XM5
timestamp 1728341492
transform 1 0 483 0 1 278
box -211 -224 211 224
<< labels >>
flabel metal1 s -150 324 -150 370 0 FreeSans 480 0 0 0 Vbias
port 4 nsew
flabel metal1 s -150 466 -150 500 0 FreeSans 480 0 0 0 Vin
port 5 nsew
flabel metal1 s -150 778 -150 812 0 FreeSans 480 0 0 0 Ctrl
port 6 nsew
flabel locali s 236 1408 308 1408 0 FreeSans 480 0 0 0 VDD
port 10 nsew
flabel locali s 236 54 308 54 0 FreeSans 480 0 0 0 GND
port 11 nsew
flabel metal1 s 694 678 694 712 0 FreeSans 480 0 0 0 Vout
port 12 nsew
<< end >>
