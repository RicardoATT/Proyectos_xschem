** sch_path: /home/ricardoatt/RATT_repos/Proyectos_xschem/opamp_design/simple_one_stage_opamp/simple_one_stage_opamp_av.sch
**.subckt simple_one_stage_opamp_av
XCL Vout VSS sky130_fd_pr__cap_mim_m3_1 W=50000000 L=1 MF=1 m=1
RL Vout VSS 100k m=1
XCL1 Vinn VSS sky130_fd_pr__cap_mim_m3_1 W=50000000 L=1 MF=1 m=1
RL1 Vout Vinn 100k m=1
V5 VDD GND 1.8
V6 Vinn GND 0.9
V7 Vinp GND ac 1 SINE(0.9 0.9 10000k)
V8 VSS GND 0
x1 VDD Vout Vinp Vinn VSS simple_one_stage_opamp
**** begin user architecture code

.ac dec 0.0001 1 1000k
.control
	run
	setplot tran1
	set color0=rgb:f/f/f
	set color1=rgb:0/0/0
	settype decibel vout
	plot vdb(Vout) xlog
	wrdata simple_one_stage_opamp_av.ssv vdb(Vout) xlog
.endc
.save all



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ricardoatt/pdk/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/ricardoatt/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ricardoatt/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ricardoatt/pdk/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/ricardoatt/RATT_repos/Proyectos_xschem/opamp_design/simple_one_stage_opamp/simple_one_stage_opamp.sym # of pins=5
** sym_path: /home/ricardoatt/RATT_repos/Proyectos_xschem/opamp_design/simple_one_stage_opamp/simple_one_stage_opamp.sym
** sch_path: /home/ricardoatt/RATT_repos/Proyectos_xschem/opamp_design/simple_one_stage_opamp/simple_one_stage_opamp.sch
.subckt simple_one_stage_opamp VDD Vout Vinp Vinn VSS
*.iopin VSS
*.iopin VDD
*.ipin Vinp
*.ipin Vinn
*.opin Vout
XM1 net2 Vinp net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=15.648 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.449 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vinn net1 VSS sky130_fd_pr__nfet_01v8 L=0.15 W=15.648 nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
XM3 Vout net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=0.449 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net1 net3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=5.193 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net3 net3 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=5.193 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I0 VDD net3 48u
.ends

.GLOBAL VDD
.GLOBAL GND
.end
