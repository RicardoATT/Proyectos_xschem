magic
tech sky130B
magscale 1 2
timestamp 1729123963
<< locali >>
rect -910 3845 -876 4027
rect -832 3998 -762 4068
rect -802 3320 -762 3460
rect -916 2996 -882 3093
rect -3424 2725 -3390 2836
rect -3016 2806 -2940 2840
rect -1870 2530 -1754 2564
rect -3424 2150 -3354 2220
rect -1724 2186 -1648 2220
rect -1536 2215 -1502 2312
rect -1242 2186 -1166 2220
<< metal1 >>
rect -3316 3923 -1008 3936
rect -3316 3890 -966 3923
rect -3316 3842 -3270 3890
rect -3124 3846 -3078 3890
rect -2932 3845 -2886 3890
rect -2740 3844 -2694 3890
rect -2548 3841 -2502 3890
rect -2356 3841 -2310 3890
rect -2164 3840 -2118 3890
rect -1972 3844 -1926 3890
rect -1780 3845 -1734 3890
rect -1588 3847 -1542 3890
rect -1396 3846 -1350 3890
rect -1204 3844 -1158 3890
rect -1012 3846 -966 3890
rect -3031 3673 -2979 3679
rect -3229 3621 -3223 3673
rect -3171 3621 -3165 3673
rect -3316 3568 -3270 3621
rect -3214 3609 -3180 3621
rect -3031 3615 -2979 3621
rect -2839 3673 -2787 3679
rect -2839 3615 -2787 3621
rect -2647 3673 -2595 3679
rect -2647 3615 -2595 3621
rect -2455 3673 -2403 3679
rect -2455 3615 -2403 3621
rect -2263 3673 -2211 3679
rect -2263 3615 -2211 3621
rect -2071 3673 -2019 3679
rect -2071 3615 -2019 3621
rect -1879 3673 -1827 3679
rect -1879 3615 -1827 3621
rect -1687 3673 -1635 3679
rect -1687 3615 -1635 3621
rect -1495 3673 -1443 3679
rect -1495 3615 -1443 3621
rect -1303 3673 -1251 3679
rect -1303 3615 -1251 3621
rect -1111 3673 -1059 3679
rect -1111 3615 -1059 3621
rect -919 3673 -867 3679
rect -919 3615 -867 3621
rect -3316 3522 -912 3568
rect -3316 3460 -3270 3522
rect -3316 3426 -3014 3460
rect -3167 3363 -3115 3369
rect -3460 3320 -3167 3354
rect -3167 3305 -3115 3311
rect -3460 3108 -3209 3142
rect -3350 2980 -3270 3070
rect -3048 3008 -3014 3426
rect -2957 3311 -2951 3363
rect -2899 3354 -2893 3363
rect -2899 3320 -2650 3354
rect -2899 3311 -2893 3320
rect -2684 3258 -2650 3320
rect -2696 3212 -1240 3258
rect -2732 3166 -2698 3168
rect -2549 3166 -2497 3172
rect -2747 3114 -2741 3166
rect -2689 3114 -2683 3166
rect -2549 3108 -2497 3114
rect -2357 3166 -2305 3172
rect -2357 3108 -2305 3114
rect -2165 3166 -2113 3172
rect -2165 3108 -2113 3114
rect -1973 3166 -1921 3172
rect -1973 3108 -1921 3114
rect -1781 3166 -1729 3172
rect -1781 3108 -1729 3114
rect -1589 3166 -1537 3172
rect -1589 3108 -1537 3114
rect -1397 3166 -1345 3172
rect -1397 3108 -1345 3114
rect -3168 2980 -2794 3008
rect -3350 2840 -3316 2980
rect -3063 2942 -3057 2951
rect -3183 2908 -3057 2942
rect -3063 2899 -3057 2908
rect -3005 2899 -2999 2951
rect -1274 2948 -1240 3212
rect -1004 3211 -912 3522
rect -2792 2902 -1240 2948
rect -2792 2840 -2730 2902
rect -3350 2806 -3276 2840
rect -3310 2749 -3276 2806
rect -3166 2806 -2730 2840
rect -2597 2849 -2545 2855
rect -3319 2743 -3267 2749
rect -3460 2700 -3390 2734
rect -3424 2220 -3390 2700
rect -3319 2685 -3267 2691
rect -3310 2546 -3276 2685
rect -3166 2638 -3132 2806
rect -1659 2849 -1607 2855
rect -2545 2806 -1659 2840
rect -2597 2791 -2545 2797
rect -1659 2791 -1607 2797
rect -2983 2743 -2931 2749
rect -2931 2700 -1259 2734
rect -2983 2685 -2931 2691
rect -1335 2652 -1259 2700
rect -3178 2592 -1722 2638
rect -1060 2630 -1014 3113
rect -966 2968 -726 3002
rect -966 2658 -932 2968
rect -3214 2550 -3180 2554
rect -3223 2544 -3171 2550
rect -3223 2486 -3171 2492
rect -3031 2544 -2979 2550
rect -3031 2486 -2979 2492
rect -2839 2544 -2787 2550
rect -2839 2486 -2787 2492
rect -2647 2544 -2595 2550
rect -2647 2486 -2595 2492
rect -2455 2544 -2403 2550
rect -2455 2486 -2403 2492
rect -2263 2544 -2211 2550
rect -2263 2486 -2211 2492
rect -2071 2544 -2019 2550
rect -2071 2486 -2019 2492
rect -1966 2487 -1932 2548
rect -1879 2544 -1827 2550
rect -1879 2486 -1827 2492
rect -3316 2424 -3270 2443
rect -3127 2424 -3075 2430
rect -3325 2372 -3319 2424
rect -3267 2372 -3261 2424
rect -3316 2366 -3270 2372
rect -3127 2366 -3075 2372
rect -2935 2424 -2883 2430
rect -2935 2366 -2883 2372
rect -2743 2424 -2691 2430
rect -2743 2366 -2691 2372
rect -2551 2424 -2499 2430
rect -2551 2366 -2499 2372
rect -2359 2424 -2307 2430
rect -2359 2366 -2307 2372
rect -2167 2424 -2115 2430
rect -2167 2366 -2115 2372
rect -1975 2424 -1923 2430
rect -1975 2366 -1923 2372
rect -1756 2328 -1722 2592
rect -1665 2519 -1659 2571
rect -1607 2519 -1601 2571
rect -1650 2460 -1616 2519
rect -1650 2426 -1416 2460
rect -1360 2385 -1323 2388
rect -1388 2339 -1323 2385
rect -1360 2336 -1323 2339
rect -1271 2336 -1265 2388
rect -3274 2282 -1722 2328
rect -1022 2220 -964 2307
rect -3424 2186 -964 2220
<< via1 >>
rect -3223 3621 -3171 3673
rect -3031 3621 -2979 3673
rect -2839 3621 -2787 3673
rect -2647 3621 -2595 3673
rect -2455 3621 -2403 3673
rect -2263 3621 -2211 3673
rect -2071 3621 -2019 3673
rect -1879 3621 -1827 3673
rect -1687 3621 -1635 3673
rect -1495 3621 -1443 3673
rect -1303 3621 -1251 3673
rect -1111 3621 -1059 3673
rect -919 3621 -867 3673
rect -3167 3311 -3115 3363
rect -2951 3311 -2899 3363
rect -2741 3114 -2689 3166
rect -2549 3114 -2497 3166
rect -2357 3114 -2305 3166
rect -2165 3114 -2113 3166
rect -1973 3114 -1921 3166
rect -1781 3114 -1729 3166
rect -1589 3114 -1537 3166
rect -1397 3114 -1345 3166
rect -3057 2899 -3005 2951
rect -3319 2691 -3267 2743
rect -2597 2797 -2545 2849
rect -1659 2797 -1607 2849
rect -2983 2691 -2931 2743
rect -3223 2492 -3171 2544
rect -3031 2492 -2979 2544
rect -2839 2492 -2787 2544
rect -2647 2492 -2595 2544
rect -2455 2492 -2403 2544
rect -2263 2492 -2211 2544
rect -2071 2492 -2019 2544
rect -1879 2492 -1827 2544
rect -3319 2372 -3267 2424
rect -3127 2372 -3075 2424
rect -2935 2372 -2883 2424
rect -2743 2372 -2691 2424
rect -2551 2372 -2499 2424
rect -2359 2372 -2307 2424
rect -2167 2372 -2115 2424
rect -1975 2372 -1923 2424
rect -1659 2519 -1607 2571
rect -1323 2336 -1271 2388
<< metal2 >>
rect -3229 3621 -3223 3673
rect -3171 3670 -3165 3673
rect -3037 3670 -3031 3673
rect -3171 3624 -3031 3670
rect -3171 3621 -3165 3624
rect -3037 3621 -3031 3624
rect -2979 3670 -2973 3673
rect -2845 3670 -2839 3673
rect -2979 3624 -2839 3670
rect -2979 3621 -2973 3624
rect -2845 3621 -2839 3624
rect -2787 3670 -2781 3673
rect -2653 3670 -2647 3673
rect -2787 3624 -2647 3670
rect -2787 3621 -2781 3624
rect -2653 3621 -2647 3624
rect -2595 3670 -2589 3673
rect -2461 3670 -2455 3673
rect -2595 3624 -2455 3670
rect -2595 3621 -2589 3624
rect -2461 3621 -2455 3624
rect -2403 3670 -2397 3673
rect -2269 3670 -2263 3673
rect -2403 3624 -2263 3670
rect -2403 3621 -2397 3624
rect -2269 3621 -2263 3624
rect -2211 3670 -2205 3673
rect -2077 3670 -2071 3673
rect -2211 3624 -2071 3670
rect -2211 3621 -2205 3624
rect -2077 3621 -2071 3624
rect -2019 3670 -2013 3673
rect -1885 3670 -1879 3673
rect -2019 3624 -1879 3670
rect -2019 3621 -2013 3624
rect -1885 3621 -1879 3624
rect -1827 3670 -1821 3673
rect -1693 3670 -1687 3673
rect -1827 3624 -1687 3670
rect -1827 3621 -1821 3624
rect -1693 3621 -1687 3624
rect -1635 3670 -1629 3673
rect -1501 3670 -1495 3673
rect -1635 3624 -1495 3670
rect -1635 3621 -1629 3624
rect -1501 3621 -1495 3624
rect -1443 3670 -1437 3673
rect -1309 3670 -1303 3673
rect -1443 3624 -1303 3670
rect -1443 3621 -1437 3624
rect -1309 3621 -1303 3624
rect -1251 3670 -1245 3673
rect -1117 3670 -1111 3673
rect -1251 3624 -1111 3670
rect -1251 3621 -1245 3624
rect -1117 3621 -1111 3624
rect -1059 3670 -1053 3673
rect -925 3670 -919 3673
rect -1059 3624 -919 3670
rect -1059 3621 -1053 3624
rect -925 3621 -919 3624
rect -867 3621 -861 3673
rect -2951 3363 -2899 3369
rect -3173 3311 -3167 3363
rect -3115 3354 -3109 3363
rect -3115 3320 -2951 3354
rect -3115 3311 -3109 3320
rect -2951 3305 -2899 3311
rect -2747 3114 -2741 3166
rect -2689 3163 -2683 3166
rect -2555 3163 -2549 3166
rect -2689 3117 -2549 3163
rect -2689 3114 -2683 3117
rect -2555 3114 -2549 3117
rect -2497 3163 -2491 3166
rect -2363 3163 -2357 3166
rect -2497 3117 -2357 3163
rect -2497 3114 -2491 3117
rect -2363 3114 -2357 3117
rect -2305 3163 -2299 3166
rect -2171 3163 -2165 3166
rect -2305 3117 -2165 3163
rect -2305 3114 -2299 3117
rect -2171 3114 -2165 3117
rect -2113 3163 -2107 3166
rect -1979 3163 -1973 3166
rect -2113 3117 -1973 3163
rect -2113 3114 -2107 3117
rect -1979 3114 -1973 3117
rect -1921 3163 -1915 3166
rect -1787 3163 -1781 3166
rect -1921 3117 -1781 3163
rect -1921 3114 -1915 3117
rect -1787 3114 -1781 3117
rect -1729 3163 -1723 3166
rect -1595 3163 -1589 3166
rect -1729 3117 -1589 3163
rect -1729 3114 -1723 3117
rect -1595 3114 -1589 3117
rect -1537 3163 -1531 3166
rect -1403 3163 -1397 3166
rect -1537 3117 -1397 3163
rect -1537 3114 -1531 3117
rect -1403 3114 -1397 3117
rect -1345 3163 -1339 3166
rect -1345 3114 -1274 3163
rect -3063 2899 -3057 2951
rect -3005 2899 -2999 2951
rect -3048 2840 -3014 2899
rect -2603 2840 -2597 2849
rect -3048 2806 -2597 2840
rect -2603 2797 -2597 2806
rect -2545 2797 -2539 2849
rect -1665 2797 -1659 2849
rect -1607 2797 -1601 2849
rect -3319 2743 -3267 2749
rect -2989 2734 -2983 2743
rect -3267 2700 -2983 2734
rect -2989 2691 -2983 2700
rect -2931 2691 -2925 2743
rect -3319 2685 -3267 2691
rect -1650 2577 -1616 2797
rect -1320 2728 -1274 3114
rect -1335 2652 -1259 2728
rect -1659 2571 -1607 2577
rect -3229 2492 -3223 2544
rect -3171 2535 -3165 2544
rect -3037 2535 -3031 2544
rect -3171 2501 -3031 2535
rect -3171 2492 -3165 2501
rect -3037 2492 -3031 2501
rect -2979 2535 -2973 2544
rect -2845 2535 -2839 2544
rect -2979 2501 -2839 2535
rect -2979 2492 -2973 2501
rect -2845 2492 -2839 2501
rect -2787 2535 -2781 2544
rect -2653 2535 -2647 2544
rect -2787 2501 -2647 2535
rect -2787 2492 -2781 2501
rect -2653 2492 -2647 2501
rect -2595 2535 -2589 2544
rect -2461 2535 -2455 2544
rect -2595 2501 -2455 2535
rect -2595 2492 -2589 2501
rect -2461 2492 -2455 2501
rect -2403 2535 -2397 2544
rect -2269 2535 -2263 2544
rect -2403 2501 -2263 2535
rect -2403 2492 -2397 2501
rect -2269 2492 -2263 2501
rect -2211 2535 -2205 2544
rect -2077 2535 -2071 2544
rect -2211 2501 -2071 2535
rect -2211 2492 -2205 2501
rect -2077 2492 -2071 2501
rect -2019 2535 -2013 2544
rect -1885 2535 -1879 2544
rect -2019 2501 -1879 2535
rect -2019 2492 -2013 2501
rect -1885 2492 -1879 2501
rect -1827 2492 -1821 2544
rect -1659 2513 -1607 2519
rect -3325 2372 -3319 2424
rect -3267 2421 -3261 2424
rect -3133 2421 -3127 2424
rect -3267 2375 -3127 2421
rect -3267 2372 -3261 2375
rect -3133 2372 -3127 2375
rect -3075 2421 -3069 2424
rect -2941 2421 -2935 2424
rect -3075 2375 -2935 2421
rect -3075 2372 -3069 2375
rect -2941 2372 -2935 2375
rect -2883 2421 -2877 2424
rect -2749 2421 -2743 2424
rect -2883 2375 -2743 2421
rect -2883 2372 -2877 2375
rect -2749 2372 -2743 2375
rect -2691 2421 -2685 2424
rect -2557 2421 -2551 2424
rect -2691 2375 -2551 2421
rect -2691 2372 -2685 2375
rect -2557 2372 -2551 2375
rect -2499 2421 -2493 2424
rect -2365 2421 -2359 2424
rect -2499 2375 -2359 2421
rect -2499 2372 -2493 2375
rect -2365 2372 -2359 2375
rect -2307 2421 -2301 2424
rect -2173 2421 -2167 2424
rect -2307 2375 -2167 2421
rect -2307 2372 -2301 2375
rect -2173 2372 -2167 2375
rect -2115 2421 -2109 2424
rect -1981 2421 -1975 2424
rect -2115 2375 -1975 2421
rect -2115 2372 -2109 2375
rect -1981 2372 -1975 2375
rect -1923 2372 -1917 2424
rect -1320 2394 -1274 2652
rect -1323 2388 -1271 2394
rect -1323 2330 -1271 2336
use sky130_fd_pr__nfet_01v8_MT8PY5  sky130_fd_pr__nfet_01v8_MT8PY5_0
timestamp 1729119800
transform 1 0 -2573 0 1 2460
box -887 -310 887 310
use sky130_fd_pr__pfet_01v8_8D7YKK  sky130_fd_pr__pfet_01v8_8D7YKK_0
timestamp 1729119800
transform 1 0 -2093 0 1 3729
box -1367 -339 1367 339
use sky130_fd_pr_reram__reram_cell  sky130_fd_pr_reram__reram_cell_0
timestamp 1727988820
transform 1 0 -1297 0 1 2690
box -38 -38 38 38
use sky130_fd_pr__nfet_01v8_KJ9A5H  XM1
timestamp 1729119800
transform -1 0 -3219 0 1 3025
box -241 -255 241 255
use sky130_fd_pr__nfet_01v8_MT8PY5  XM3
timestamp 1729119800
transform 1 0 -2091 0 1 3080
box -887 -310 887 310
use sky130_fd_pr__nfet_01v8_P46M8Q  XM4
timestamp 1729119800
transform -1 0 -1445 0 1 2374
box -241 -224 241 224
use sky130_fd_pr__pfet_01v8_5M8GQ7  XM6
timestamp 1729119800
transform 1 0 -968 0 1 3161
box -236 -229 236 229
use sky130_fd_pr__nfet_01v8_84QSGM  XM7
timestamp 1729119800
transform 1 0 -993 0 1 2479
box -211 -329 211 329
<< labels >>
flabel metal1 s -726 2968 -726 3002 0 FreeSans 480 0 0 0 Ipos
port 24 nsew
flabel metal1 s -3460 3320 -3460 3354 0 FreeSans 480 0 0 0 Vpos
port 25 nsew
flabel metal1 s -3460 3108 -3460 3142 0 FreeSans 480 0 0 0 Vpre
port 26 nsew
flabel metal1 s -3460 2700 -3460 2734 0 FreeSans 480 0 0 0 ctrl_pos
port 27 nsew
flabel locali s -3424 2150 -3354 2150 0 FreeSans 480 0 0 0 GND
port 28 nsew
flabel locali s -832 4068 -762 4068 0 FreeSans 480 0 0 0 VDD
port 29 nsew
<< end >>
