* SPICE3 file created from Syn_7T1R.ext - technology: sky130B

.subckt Syn_7T1R Vpos ctrl_pos Vpre Ipos GND VDD
C0 XM6/G sky130_fd_pr__nfet_01v8_X2WNKZ_0/S 2.427512f
C1 XM6/G VDD 6.266848f
Xsky130_fd_pr__nfet_01v8_P46M8Q_0 Vpre sky130_fd_pr__nfet_01v8_X2WNKZ_0/S GND GND
+ sky130_fd_pr__nfet_01v8_P46M8Q
Xsky130_fd_pr_reram__reram_cell_0 sky130_fd_pr__nfet_01v8_X2WNKZ_0/S XM2/D sky130_fd_pr_reram__reram_cell
XXM1 Vpre XM6/G XM2/D GND sky130_fd_pr__nfet_01v8_P46M8Q
XXM2 Vpos XM2/D GND GND sky130_fd_pr__nfet_01v8_X2WNKZ
XXM5 XM6/G XM6/G VDD VDD sky130_fd_pr__pfet_01v8_UGKMGH
XXM6 VDD XM6/G XM7/D VDD sky130_fd_pr__pfet_01v8_UAJFQ5
XXM7 ctrl_pos XM7/D Ipos GND sky130_fd_pr__nfet_01v8_84QSGM
Xsky130_fd_pr__nfet_01v8_X2WNKZ_0 Vpos XM6/G sky130_fd_pr__nfet_01v8_X2WNKZ_0/S GND
+ sky130_fd_pr__nfet_01v8_X2WNKZ
C2 VDD GND 7.550229f
C3 XM6/G GND 2.418188f
C4 XM2/D GND 3.94803f
C5 Vpre GND 2.643731f
.ends
