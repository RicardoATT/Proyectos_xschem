magic
tech sky130B
magscale 1 2
timestamp 1728435493
<< error_p >>
rect -29 -157 29 -151
rect -29 -191 -17 -157
rect -29 -197 29 -191
<< pwell >>
rect -211 -329 211 329
<< nmos >>
rect -15 -119 15 181
<< ndiff >>
rect -73 169 -15 181
rect -73 -107 -61 169
rect -27 -107 -15 169
rect -73 -119 -15 -107
rect 15 169 73 181
rect 15 -107 27 169
rect 61 -107 73 169
rect 15 -119 73 -107
<< ndiffc >>
rect -61 -107 -27 169
rect 27 -107 61 169
<< psubdiff >>
rect -175 259 -79 293
rect 79 259 175 293
rect -175 197 -141 259
rect 141 197 175 259
rect -175 -259 -141 -197
rect 141 -259 175 -197
rect -175 -293 -79 -259
rect 79 -293 175 -259
<< psubdiffcont >>
rect -79 259 79 293
rect -175 -197 -141 197
rect 141 -197 175 197
rect -79 -293 79 -259
<< poly >>
rect -15 181 15 207
rect -15 -141 15 -119
rect -33 -157 33 -141
rect -33 -191 -17 -157
rect 17 -191 33 -157
rect -33 -207 33 -191
<< polycont >>
rect -17 -191 17 -157
<< locali >>
rect -175 259 -79 293
rect 79 259 175 293
rect -175 197 -141 259
rect 141 197 175 259
rect -61 169 -27 185
rect -61 -123 -27 -107
rect 27 169 61 185
rect 27 -123 61 -107
rect -33 -191 -17 -157
rect 17 -191 33 -157
rect -175 -259 -141 -197
rect 141 -259 175 -197
rect -175 -293 -79 -259
rect 79 -293 175 -259
<< viali >>
rect -61 -107 -27 169
rect 27 -107 61 169
rect -17 -191 17 -157
<< metal1 >>
rect -67 169 -21 181
rect -67 -107 -61 169
rect -27 -107 -21 169
rect -67 -119 -21 -107
rect 21 169 67 181
rect 21 -107 27 169
rect 61 -107 67 169
rect 21 -119 67 -107
rect -29 -157 29 -151
rect -29 -191 -17 -157
rect 17 -191 29 -157
rect -29 -197 29 -191
<< labels >>
flabel metal1 s 0 -174 0 -174 0 FreeSans 480 0 0 0 G
port 8 nsew
flabel metal1 s -44 32 -44 32 0 FreeSans 480 0 0 0 D
port 9 nsew
flabel metal1 s 44 30 44 30 0 FreeSans 480 0 0 0 S
port 10 nsew
flabel locali s 0 -275 0 -275 0 FreeSans 480 0 0 0 B
port 11 nsew
<< properties >>
string FIXED_BBOX -158 -276 158 276
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
