magic
tech sky130B
magscale 1 2
timestamp 1729119800
<< pwell >>
rect -241 -255 241 255
<< nmos >>
rect -45 -45 45 45
<< ndiff >>
rect -103 33 -45 45
rect -103 -33 -91 33
rect -57 -33 -45 33
rect -103 -45 -45 -33
rect 45 33 103 45
rect 45 -33 57 33
rect 91 -33 103 33
rect 45 -45 103 -33
<< ndiffc >>
rect -91 -33 -57 33
rect 57 -33 91 33
<< psubdiff >>
rect -205 185 -109 219
rect 109 185 205 219
rect -205 123 -171 185
rect 171 123 205 185
rect -205 -185 -171 -123
rect 171 -185 205 -123
rect -205 -219 -109 -185
rect 109 -219 205 -185
<< psubdiffcont >>
rect -109 185 109 219
rect -205 -123 -171 123
rect 171 -123 205 123
rect -109 -219 109 -185
<< poly >>
rect -45 117 45 133
rect -45 83 -29 117
rect 29 83 45 117
rect -45 45 45 83
rect -45 -83 45 -45
rect -45 -117 -29 -83
rect 29 -117 45 -83
rect -45 -133 45 -117
<< polycont >>
rect -29 83 29 117
rect -29 -117 29 -83
<< locali >>
rect -205 185 -109 219
rect 109 185 205 219
rect -205 123 -171 185
rect 171 123 205 185
rect -45 83 -29 117
rect 29 83 45 117
rect -91 33 -57 49
rect -91 -49 -57 -33
rect 57 33 91 49
rect 57 -49 91 -33
rect -45 -117 -29 -83
rect 29 -117 45 -83
rect -205 -185 -171 -123
rect 171 -185 205 -123
rect -205 -219 -109 -185
rect 109 -219 205 -185
<< viali >>
rect -29 83 29 117
rect -91 -33 -57 33
rect 57 -33 91 33
rect -29 -117 29 -83
<< metal1 >>
rect -41 117 41 123
rect -41 83 -29 117
rect 29 83 41 117
rect -41 77 41 83
rect -97 33 -51 45
rect -97 -33 -91 33
rect -57 -33 -51 33
rect -97 -45 -51 -33
rect 51 33 97 45
rect 51 -33 57 33
rect 91 -33 97 33
rect 51 -45 97 -33
rect -41 -83 41 -77
rect -41 -117 -29 -83
rect 29 -117 41 -83
rect -41 -123 41 -117
<< labels >>
flabel locali s 0 201 0 201 0 FreeSans 480 0 0 0 B
port 4 nsew
flabel metal1 s 2 99 2 99 0 FreeSans 480 0 0 0 G
port 5 nsew
flabel metal1 s -74 -1 -74 -1 0 FreeSans 480 0 0 0 D
port 6 nsew
flabel metal1 s 75 -2 75 -2 0 FreeSans 480 0 0 0 S
port 7 nsew
<< properties >>
string FIXED_BBOX -188 -202 188 202
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 0.45 l 0.45 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
