** sch_path: /home/ricardo/RATT-repo/Proyectos-RATT/Proyectos-xschem/inverter/inverter_tb.sch
**.subckt inverter_tb
x1 net1 vout vin GND inverter
V1 vin GND PULSE(0 1.8 0 1n 1n 50n 100n 4)
.save i(v1)
V2 net1 GND 1.8
.save i(v2)
**** begin user architecture code


.control
	save all
	run
	tran 10p 400n
	write inverter_tb.raw
.endc



** opencircuitdesign pdks install
.lib /home/ricardo/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt


**** end user architecture code
**.ends

* expanding   symbol:  /home/ricardo/Escritorio/Proyectos_xschem/inverter/inverter.sym # of pins=4
** sym_path: /home/ricardo/Escritorio/Proyectos_xschem/inverter/inverter.sym
** sch_path: /home/ricardo/Escritorio/Proyectos_xschem/inverter/inverter.sch
.subckt inverter vdd vout vin gnd
*.ipin vin
*.iopin vdd
*.opin vout
*.iopin gnd
XM1 vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 vout vin gnd gnd sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.GLOBAL GND
.end
