magic
tech sky130B
magscale 1 2
timestamp 1728505772
<< locali >>
rect -689 6185 -619 6255
rect -803 5753 -769 5840
rect -971 5437 -857 5471
rect -689 -525 -655 6185
rect -583 5480 -549 6218
rect -469 5757 -435 5844
rect -583 5446 -435 5480
rect -583 4912 -549 5446
rect -583 4878 -435 4912
rect -583 4344 -549 4878
rect -583 4310 -435 4344
rect -583 3776 -549 4310
rect -583 3742 -435 3776
rect -583 3208 -549 3742
rect -583 3174 -435 3208
rect -583 2640 -549 3174
rect -583 2606 -435 2640
rect -583 2072 -549 2606
rect -583 2038 -435 2072
rect -583 1504 -549 2038
rect -583 1470 -435 1504
rect -583 936 -549 1470
rect -583 902 -435 936
rect -583 368 -549 902
rect -583 334 -435 368
rect -583 -200 -549 334
rect -583 -234 -435 -200
rect -583 -482 -549 -234
rect -619 -561 -549 -482
<< metal1 >>
rect -937 6218 -903 6219
rect -937 6185 -301 6218
rect -937 6035 -903 6185
rect -847 6082 -391 6116
rect -937 6007 -857 6035
rect -1041 5617 -813 5651
rect -847 5548 -813 5617
rect -583 5650 -549 6082
rect -335 6044 -301 6185
rect -381 6016 -233 6044
rect -583 5616 -301 5650
rect -847 5514 -391 5548
rect -335 5476 -301 5616
rect -381 5448 -301 5476
rect -698 5307 -646 5313
rect -763 5267 -698 5295
rect -381 5276 -301 5304
rect -698 5249 -646 5255
rect -1041 5049 -813 5083
rect -847 4980 -813 5049
rect -847 4946 -391 4980
rect -704 4899 -698 4912
rect -763 4871 -698 4899
rect -704 4860 -698 4871
rect -646 4860 -640 4912
rect -335 4908 -301 5276
rect -381 4880 -301 4908
rect -937 4699 -897 4727
rect -381 4708 -301 4736
rect -1017 4524 -965 4530
rect -1041 4481 -1017 4515
rect -1017 4466 -965 4472
rect -937 4331 -903 4699
rect -856 4524 -804 4530
rect -856 4466 -804 4472
rect -847 4412 -813 4466
rect -847 4378 -391 4412
rect -335 4340 -301 4708
rect -937 4303 -897 4331
rect -381 4312 -301 4340
rect -698 4171 -646 4177
rect -763 4131 -698 4159
rect -381 4140 -301 4168
rect -698 4113 -646 4119
rect -1041 3913 -813 3947
rect -847 3844 -813 3913
rect -847 3810 -391 3844
rect -704 3763 -698 3775
rect -763 3735 -698 3763
rect -704 3723 -698 3735
rect -646 3723 -640 3775
rect -335 3772 -301 4140
rect -381 3744 -301 3772
rect -937 3563 -897 3591
rect -381 3572 -301 3600
rect -1017 3388 -965 3394
rect -1041 3345 -1017 3379
rect -1017 3330 -965 3336
rect -937 3195 -903 3563
rect -856 3388 -804 3394
rect -856 3330 -804 3336
rect -847 3276 -813 3330
rect -847 3242 -391 3276
rect -335 3204 -301 3572
rect -937 3167 -897 3195
rect -381 3176 -301 3204
rect -704 3023 -698 3035
rect -763 2995 -698 3023
rect -704 2983 -698 2995
rect -646 2983 -640 3035
rect -381 3004 -301 3032
rect -1041 2777 -813 2811
rect -847 2708 -813 2777
rect -847 2674 -391 2708
rect -704 2627 -698 2639
rect -763 2599 -698 2627
rect -704 2587 -698 2599
rect -646 2587 -640 2639
rect -335 2636 -301 3004
rect -267 2868 -233 6016
rect -267 2834 -197 2868
rect -381 2608 -301 2636
rect -937 2427 -897 2455
rect -381 2436 -301 2464
rect -1017 2252 -965 2258
rect -1041 2209 -1017 2243
rect -1017 2194 -965 2200
rect -937 2059 -903 2427
rect -856 2252 -804 2258
rect -856 2194 -804 2200
rect -847 2140 -813 2194
rect -847 2106 -391 2140
rect -335 2068 -301 2436
rect -937 2031 -897 2059
rect -381 2040 -301 2068
rect -704 1887 -698 1899
rect -763 1859 -698 1887
rect -704 1847 -698 1859
rect -646 1847 -640 1899
rect -381 1868 -301 1896
rect -1041 1641 -813 1675
rect -847 1572 -813 1641
rect -847 1538 -391 1572
rect -704 1491 -698 1503
rect -763 1463 -698 1491
rect -704 1451 -698 1463
rect -646 1451 -640 1503
rect -335 1500 -301 1868
rect -381 1472 -301 1500
rect -937 1291 -897 1319
rect -381 1300 -301 1328
rect -1017 1116 -965 1122
rect -1041 1073 -1017 1107
rect -1017 1058 -965 1064
rect -937 923 -903 1291
rect -856 1116 -804 1122
rect -856 1058 -804 1064
rect -847 1004 -813 1058
rect -847 970 -391 1004
rect -335 932 -301 1300
rect -937 895 -897 923
rect -381 904 -301 932
rect -704 751 -698 763
rect -763 723 -698 751
rect -704 711 -698 723
rect -646 711 -640 763
rect -381 732 -301 760
rect -1041 505 -813 539
rect -847 430 -813 505
rect -847 396 -391 430
rect -704 355 -698 367
rect -763 327 -698 355
rect -704 315 -698 327
rect -646 315 -640 367
rect -335 364 -301 732
rect -381 336 -301 364
rect -937 155 -897 183
rect -381 164 -301 192
rect -1017 -20 -965 -14
rect -1041 -63 -1017 -29
rect -1017 -78 -965 -72
rect -937 -213 -903 155
rect -856 -20 -804 -14
rect -856 -78 -804 -72
rect -847 -138 -813 -78
rect -847 -172 -391 -138
rect -335 -204 -301 164
rect -937 -241 -897 -213
rect -381 -232 -301 -204
rect -381 -404 -341 -376
<< via1 >>
rect -698 5255 -646 5307
rect -698 4860 -646 4912
rect -1017 4472 -965 4524
rect -856 4472 -804 4524
rect -698 4119 -646 4171
rect -698 3723 -646 3775
rect -1017 3336 -965 3388
rect -856 3336 -804 3388
rect -698 2983 -646 3035
rect -698 2587 -646 2639
rect -1017 2200 -965 2252
rect -856 2200 -804 2252
rect -698 1847 -646 1899
rect -698 1451 -646 1503
rect -1017 1064 -965 1116
rect -856 1064 -804 1116
rect -698 711 -646 763
rect -698 315 -646 367
rect -1017 -72 -965 -20
rect -856 -72 -804 -20
<< metal2 >>
rect -704 5255 -698 5307
rect -646 5255 -640 5307
rect -689 4918 -655 5255
rect -698 4912 -646 4918
rect -698 4854 -646 4860
rect -1023 4472 -1017 4524
rect -965 4515 -959 4524
rect -862 4515 -856 4524
rect -965 4481 -856 4515
rect -965 4472 -959 4481
rect -862 4472 -856 4481
rect -804 4472 -798 4524
rect -704 4119 -698 4171
rect -646 4119 -640 4171
rect -689 3781 -655 4119
rect -698 3775 -646 3781
rect -698 3717 -646 3723
rect -1023 3336 -1017 3388
rect -965 3379 -959 3388
rect -862 3379 -856 3388
rect -965 3345 -856 3379
rect -965 3336 -959 3345
rect -862 3336 -856 3345
rect -804 3336 -798 3388
rect -698 3035 -646 3041
rect -698 2977 -646 2983
rect -689 2645 -655 2977
rect -698 2639 -646 2645
rect -698 2581 -646 2587
rect -1023 2200 -1017 2252
rect -965 2243 -959 2252
rect -862 2243 -856 2252
rect -965 2209 -856 2243
rect -965 2200 -959 2209
rect -862 2200 -856 2209
rect -804 2200 -798 2252
rect -698 1899 -646 1905
rect -698 1841 -646 1847
rect -689 1509 -655 1841
rect -698 1503 -646 1509
rect -698 1445 -646 1451
rect -1023 1064 -1017 1116
rect -965 1107 -959 1116
rect -862 1107 -856 1116
rect -965 1073 -856 1107
rect -965 1064 -959 1073
rect -862 1064 -856 1073
rect -804 1064 -798 1116
rect -698 763 -646 769
rect -698 705 -646 711
rect -689 373 -655 705
rect -698 367 -646 373
rect -698 309 -646 315
rect -1023 -72 -1017 -20
rect -965 -29 -959 -20
rect -862 -29 -856 -20
rect -965 -63 -856 -29
rect -965 -72 -959 -63
rect -862 -72 -856 -63
rect -804 -72 -798 -20
use sky130_fd_pr__nfet_01v8_64Z3AY  sky130_fd_pr__nfet_01v8_64Z3AY_0
timestamp 1728500067
transform 1 0 -408 0 1 5407
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  sky130_fd_pr__pfet_01v8_MGS3BN_0
timestamp 1728412239
transform 1 0 -830 0 1 5403
box -211 -284 211 284
use sky130_fd_pr__pfet_01v8_MGS3BN  XM1
timestamp 1728412239
transform -1 0 -830 0 1 5971
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1728500067
transform 1 0 -408 0 1 5975
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM3
timestamp 1728412239
transform 1 0 -830 0 1 -277
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM4
timestamp 1728500067
transform 1 0 -408 0 1 -273
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM5
timestamp 1728412239
transform -1 0 -830 0 1 291
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM6
timestamp 1728500067
transform 1 0 -408 0 1 295
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM7
timestamp 1728412239
transform 1 0 -830 0 1 859
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM8
timestamp 1728500067
transform 1 0 -408 0 1 863
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM9
timestamp 1728412239
transform -1 0 -830 0 1 1427
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM10
timestamp 1728500067
transform 1 0 -408 0 1 1431
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM11
timestamp 1728412239
transform 1 0 -830 0 1 1995
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM12
timestamp 1728500067
transform 1 0 -408 0 1 1999
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM13
timestamp 1728412239
transform -1 0 -830 0 1 2563
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM14
timestamp 1728500067
transform 1 0 -408 0 1 2567
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM15
timestamp 1728412239
transform 1 0 -830 0 1 3131
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM16
timestamp 1728500067
transform 1 0 -408 0 1 3135
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM17
timestamp 1728412239
transform -1 0 -830 0 1 3699
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM18
timestamp 1728500067
transform 1 0 -408 0 1 3703
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM19
timestamp 1728412239
transform 1 0 -830 0 1 4267
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM20
timestamp 1728500067
transform 1 0 -408 0 1 4271
box -211 -279 211 279
use sky130_fd_pr__pfet_01v8_MGS3BN  XM21
timestamp 1728412239
transform -1 0 -830 0 1 4835
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM22
timestamp 1728500067
transform 1 0 -408 0 1 4839
box -211 -279 211 279
<< labels >>
flabel metal1 s -197 2834 -197 2868 0 FreeSans 480 0 0 0 out
port 0 nsew
flabel metal1 s -1041 -63 -1041 -29 0 FreeSans 480 0 0 0 N0
port 1 nsew
flabel metal1 s -1041 505 -1041 539 0 FreeSans 480 0 0 0 N1
port 2 nsew
flabel metal1 s -1041 1073 -1041 1107 0 FreeSans 480 0 0 0 N2
port 3 nsew
flabel metal1 s -1041 1641 -1041 1675 0 FreeSans 480 0 0 0 N3
port 4 nsew
flabel metal1 s -1041 2209 -1041 2243 0 FreeSans 480 0 0 0 N4
port 5 nsew
flabel metal1 s -1041 2777 -1041 2811 0 FreeSans 480 0 0 0 N5
port 6 nsew
flabel metal1 s -1041 3345 -1041 3379 0 FreeSans 480 0 0 0 N6
port 7 nsew
flabel metal1 s -1041 3913 -1041 3947 0 FreeSans 480 0 0 0 N7
port 8 nsew
flabel metal1 s -1041 4481 -1041 4515 0 FreeSans 480 0 0 0 N8
port 9 nsew
flabel metal1 s -1041 5049 -1041 5083 0 FreeSans 480 0 0 0 N9
port 10 nsew
flabel metal1 s -1041 5617 -1041 5651 0 FreeSans 480 0 0 0 RST
port 11 nsew
flabel locali s -689 6255 -619 6255 0 FreeSans 480 0 0 0 vdd
port 12 nsew
flabel locali s -619 -561 -549 -561 0 FreeSans 480 0 0 0 gnd
port 13 nsew
<< end >>
