magic
tech sky130B
magscale 1 2
timestamp 1728435493
<< error_p >>
rect -36 -56 36 -50
rect -36 -90 -24 -56
rect -36 -96 36 -90
<< nwell >>
rect -236 -229 236 229
<< pmos >>
rect -40 -9 40 81
<< pdiff >>
rect -98 69 -40 81
rect -98 3 -86 69
rect -52 3 -40 69
rect -98 -9 -40 3
rect 40 69 98 81
rect 40 3 52 69
rect 86 3 98 69
rect 40 -9 98 3
<< pdiffc >>
rect -86 3 -52 69
rect 52 3 86 69
<< nsubdiff >>
rect -200 159 -104 193
rect 104 159 200 193
rect -200 96 -166 159
rect 166 96 200 159
rect -200 -159 -166 -96
rect 166 -159 200 -96
rect -200 -193 -104 -159
rect 104 -193 200 -159
<< nsubdiffcont >>
rect -104 159 104 193
rect -200 -96 -166 96
rect 166 -96 200 96
rect -104 -193 104 -159
<< poly >>
rect -40 81 40 107
rect -40 -56 40 -9
rect -40 -90 -24 -56
rect 24 -90 40 -56
rect -40 -106 40 -90
<< polycont >>
rect -24 -90 24 -56
<< locali >>
rect -200 159 -104 193
rect 104 159 200 193
rect -200 96 -166 159
rect 166 96 200 159
rect -86 69 -52 85
rect -86 -13 -52 3
rect 52 69 86 85
rect 52 -13 86 3
rect -40 -90 -24 -56
rect 24 -90 40 -56
rect -200 -159 -166 -96
rect 166 -159 200 -96
rect -200 -193 -104 -159
rect 104 -193 200 -159
<< viali >>
rect -86 3 -52 69
rect 52 3 86 69
rect -24 -90 24 -56
<< metal1 >>
rect -92 69 -46 81
rect -92 3 -86 69
rect -52 3 -46 69
rect -92 -9 -46 3
rect 46 69 92 81
rect 46 3 52 69
rect 86 3 92 69
rect 46 -9 92 3
rect -36 -56 36 -50
rect -36 -90 -24 -56
rect 24 -90 36 -56
rect -36 -96 36 -90
<< labels >>
flabel locali s 0 176 0 176 0 FreeSans 480 0 0 0 B
port 12 nsew
flabel metal1 s 0 -73 0 -73 0 FreeSans 480 0 0 0 G
port 13 nsew
flabel metal1 s -69 35 -69 35 0 FreeSans 480 0 0 0 D
port 14 nsew
flabel metal1 s 69 34 69 34 0 FreeSans 480 0 0 0 S
port 15 nsew
<< properties >>
string FIXED_BBOX -183 -176 183 176
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.45 l 0.4 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
