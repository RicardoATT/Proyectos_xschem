magic
tech sky130B
magscale 1 2
timestamp 1729119800
<< error_p >>
rect -1325 181 -1267 187
rect -1133 181 -1075 187
rect -941 181 -883 187
rect -749 181 -691 187
rect -557 181 -499 187
rect -365 181 -307 187
rect -173 181 -115 187
rect 19 181 77 187
rect 211 181 269 187
rect 403 181 461 187
rect 595 181 653 187
rect 787 181 845 187
rect 979 181 1037 187
rect 1171 181 1229 187
rect 1363 181 1421 187
rect -1325 147 -1313 181
rect -1133 147 -1121 181
rect -941 147 -929 181
rect -749 147 -737 181
rect -557 147 -545 181
rect -365 147 -353 181
rect -173 147 -161 181
rect 19 147 31 181
rect 211 147 223 181
rect 403 147 415 181
rect 595 147 607 181
rect 787 147 799 181
rect 979 147 991 181
rect 1171 147 1183 181
rect 1363 147 1375 181
rect -1325 141 -1267 147
rect -1133 141 -1075 147
rect -941 141 -883 147
rect -749 141 -691 147
rect -557 141 -499 147
rect -365 141 -307 147
rect -173 141 -115 147
rect 19 141 77 147
rect 211 141 269 147
rect 403 141 461 147
rect 595 141 653 147
rect 787 141 845 147
rect 979 141 1037 147
rect 1171 141 1229 147
rect 1363 141 1421 147
rect -1421 -147 -1363 -141
rect -1229 -147 -1171 -141
rect -1037 -147 -979 -141
rect -845 -147 -787 -141
rect -653 -147 -595 -141
rect -461 -147 -403 -141
rect -269 -147 -211 -141
rect -77 -147 -19 -141
rect 115 -147 173 -141
rect 307 -147 365 -141
rect 499 -147 557 -141
rect 691 -147 749 -141
rect 883 -147 941 -141
rect 1075 -147 1133 -141
rect 1267 -147 1325 -141
rect -1421 -181 -1409 -147
rect -1229 -181 -1217 -147
rect -1037 -181 -1025 -147
rect -845 -181 -833 -147
rect -653 -181 -641 -147
rect -461 -181 -449 -147
rect -269 -181 -257 -147
rect -77 -181 -65 -147
rect 115 -181 127 -147
rect 307 -181 319 -147
rect 499 -181 511 -147
rect 691 -181 703 -147
rect 883 -181 895 -147
rect 1075 -181 1087 -147
rect 1267 -181 1279 -147
rect -1421 -187 -1363 -181
rect -1229 -187 -1171 -181
rect -1037 -187 -979 -181
rect -845 -187 -787 -181
rect -653 -187 -595 -181
rect -461 -187 -403 -181
rect -269 -187 -211 -181
rect -77 -187 -19 -181
rect 115 -187 173 -181
rect 307 -187 365 -181
rect 499 -187 557 -181
rect 691 -187 749 -181
rect 883 -187 941 -181
rect 1075 -187 1133 -181
rect 1267 -187 1325 -181
<< nwell >>
rect -1607 -319 1607 319
<< pmos >>
rect -1407 -100 -1377 100
rect -1311 -100 -1281 100
rect -1215 -100 -1185 100
rect -1119 -100 -1089 100
rect -1023 -100 -993 100
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
rect 993 -100 1023 100
rect 1089 -100 1119 100
rect 1185 -100 1215 100
rect 1281 -100 1311 100
rect 1377 -100 1407 100
<< pdiff >>
rect -1469 88 -1407 100
rect -1469 -88 -1457 88
rect -1423 -88 -1407 88
rect -1469 -100 -1407 -88
rect -1377 88 -1311 100
rect -1377 -88 -1361 88
rect -1327 -88 -1311 88
rect -1377 -100 -1311 -88
rect -1281 88 -1215 100
rect -1281 -88 -1265 88
rect -1231 -88 -1215 88
rect -1281 -100 -1215 -88
rect -1185 88 -1119 100
rect -1185 -88 -1169 88
rect -1135 -88 -1119 88
rect -1185 -100 -1119 -88
rect -1089 88 -1023 100
rect -1089 -88 -1073 88
rect -1039 -88 -1023 88
rect -1089 -100 -1023 -88
rect -993 88 -927 100
rect -993 -88 -977 88
rect -943 -88 -927 88
rect -993 -100 -927 -88
rect -897 88 -831 100
rect -897 -88 -881 88
rect -847 -88 -831 88
rect -897 -100 -831 -88
rect -801 88 -735 100
rect -801 -88 -785 88
rect -751 -88 -735 88
rect -801 -100 -735 -88
rect -705 88 -639 100
rect -705 -88 -689 88
rect -655 -88 -639 88
rect -705 -100 -639 -88
rect -609 88 -543 100
rect -609 -88 -593 88
rect -559 -88 -543 88
rect -609 -100 -543 -88
rect -513 88 -447 100
rect -513 -88 -497 88
rect -463 -88 -447 88
rect -513 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 513 100
rect 447 -88 463 88
rect 497 -88 513 88
rect 447 -100 513 -88
rect 543 88 609 100
rect 543 -88 559 88
rect 593 -88 609 88
rect 543 -100 609 -88
rect 639 88 705 100
rect 639 -88 655 88
rect 689 -88 705 88
rect 639 -100 705 -88
rect 735 88 801 100
rect 735 -88 751 88
rect 785 -88 801 88
rect 735 -100 801 -88
rect 831 88 897 100
rect 831 -88 847 88
rect 881 -88 897 88
rect 831 -100 897 -88
rect 927 88 993 100
rect 927 -88 943 88
rect 977 -88 993 88
rect 927 -100 993 -88
rect 1023 88 1089 100
rect 1023 -88 1039 88
rect 1073 -88 1089 88
rect 1023 -100 1089 -88
rect 1119 88 1185 100
rect 1119 -88 1135 88
rect 1169 -88 1185 88
rect 1119 -100 1185 -88
rect 1215 88 1281 100
rect 1215 -88 1231 88
rect 1265 -88 1281 88
rect 1215 -100 1281 -88
rect 1311 88 1377 100
rect 1311 -88 1327 88
rect 1361 -88 1377 88
rect 1311 -100 1377 -88
rect 1407 88 1469 100
rect 1407 -88 1423 88
rect 1457 -88 1469 88
rect 1407 -100 1469 -88
<< pdiffc >>
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
<< nsubdiff >>
rect -1571 249 -1475 283
rect 1475 249 1571 283
rect -1571 187 -1537 249
rect 1537 187 1571 249
rect -1571 -249 -1537 -187
rect 1537 -249 1571 -187
rect -1571 -283 -1475 -249
rect 1475 -283 1571 -249
<< nsubdiffcont >>
rect -1475 249 1475 283
rect -1571 -187 -1537 187
rect 1537 -187 1571 187
rect -1475 -283 1475 -249
<< poly >>
rect -1329 181 -1263 197
rect -1329 147 -1313 181
rect -1279 147 -1263 181
rect -1329 131 -1263 147
rect -1137 181 -1071 197
rect -1137 147 -1121 181
rect -1087 147 -1071 181
rect -1137 131 -1071 147
rect -945 181 -879 197
rect -945 147 -929 181
rect -895 147 -879 181
rect -945 131 -879 147
rect -753 181 -687 197
rect -753 147 -737 181
rect -703 147 -687 181
rect -753 131 -687 147
rect -561 181 -495 197
rect -561 147 -545 181
rect -511 147 -495 181
rect -561 131 -495 147
rect -369 181 -303 197
rect -369 147 -353 181
rect -319 147 -303 181
rect -369 131 -303 147
rect -177 181 -111 197
rect -177 147 -161 181
rect -127 147 -111 181
rect -177 131 -111 147
rect 15 181 81 197
rect 15 147 31 181
rect 65 147 81 181
rect 15 131 81 147
rect 207 181 273 197
rect 207 147 223 181
rect 257 147 273 181
rect 207 131 273 147
rect 399 181 465 197
rect 399 147 415 181
rect 449 147 465 181
rect 399 131 465 147
rect 591 181 657 197
rect 591 147 607 181
rect 641 147 657 181
rect 591 131 657 147
rect 783 181 849 197
rect 783 147 799 181
rect 833 147 849 181
rect 783 131 849 147
rect 975 181 1041 197
rect 975 147 991 181
rect 1025 147 1041 181
rect 975 131 1041 147
rect 1167 181 1233 197
rect 1167 147 1183 181
rect 1217 147 1233 181
rect 1167 131 1233 147
rect 1359 181 1425 197
rect 1359 147 1375 181
rect 1409 147 1425 181
rect 1359 131 1425 147
rect -1407 100 -1377 126
rect -1311 100 -1281 131
rect -1215 100 -1185 126
rect -1119 100 -1089 131
rect -1023 100 -993 126
rect -927 100 -897 131
rect -831 100 -801 126
rect -735 100 -705 131
rect -639 100 -609 126
rect -543 100 -513 131
rect -447 100 -417 126
rect -351 100 -321 131
rect -255 100 -225 126
rect -159 100 -129 131
rect -63 100 -33 126
rect 33 100 63 131
rect 129 100 159 126
rect 225 100 255 131
rect 321 100 351 126
rect 417 100 447 131
rect 513 100 543 126
rect 609 100 639 131
rect 705 100 735 126
rect 801 100 831 131
rect 897 100 927 126
rect 993 100 1023 131
rect 1089 100 1119 126
rect 1185 100 1215 131
rect 1281 100 1311 126
rect 1377 100 1407 131
rect -1407 -131 -1377 -100
rect -1311 -126 -1281 -100
rect -1215 -131 -1185 -100
rect -1119 -126 -1089 -100
rect -1023 -131 -993 -100
rect -927 -126 -897 -100
rect -831 -131 -801 -100
rect -735 -126 -705 -100
rect -639 -131 -609 -100
rect -543 -126 -513 -100
rect -447 -131 -417 -100
rect -351 -126 -321 -100
rect -255 -131 -225 -100
rect -159 -126 -129 -100
rect -63 -131 -33 -100
rect 33 -126 63 -100
rect 129 -131 159 -100
rect 225 -126 255 -100
rect 321 -131 351 -100
rect 417 -126 447 -100
rect 513 -131 543 -100
rect 609 -126 639 -100
rect 705 -131 735 -100
rect 801 -126 831 -100
rect 897 -131 927 -100
rect 993 -126 1023 -100
rect 1089 -131 1119 -100
rect 1185 -126 1215 -100
rect 1281 -131 1311 -100
rect 1377 -126 1407 -100
rect -1425 -147 -1359 -131
rect -1425 -181 -1409 -147
rect -1375 -181 -1359 -147
rect -1425 -197 -1359 -181
rect -1233 -147 -1167 -131
rect -1233 -181 -1217 -147
rect -1183 -181 -1167 -147
rect -1233 -197 -1167 -181
rect -1041 -147 -975 -131
rect -1041 -181 -1025 -147
rect -991 -181 -975 -147
rect -1041 -197 -975 -181
rect -849 -147 -783 -131
rect -849 -181 -833 -147
rect -799 -181 -783 -147
rect -849 -197 -783 -181
rect -657 -147 -591 -131
rect -657 -181 -641 -147
rect -607 -181 -591 -147
rect -657 -197 -591 -181
rect -465 -147 -399 -131
rect -465 -181 -449 -147
rect -415 -181 -399 -147
rect -465 -197 -399 -181
rect -273 -147 -207 -131
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -273 -197 -207 -181
rect -81 -147 -15 -131
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect -81 -197 -15 -181
rect 111 -147 177 -131
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 111 -197 177 -181
rect 303 -147 369 -131
rect 303 -181 319 -147
rect 353 -181 369 -147
rect 303 -197 369 -181
rect 495 -147 561 -131
rect 495 -181 511 -147
rect 545 -181 561 -147
rect 495 -197 561 -181
rect 687 -147 753 -131
rect 687 -181 703 -147
rect 737 -181 753 -147
rect 687 -197 753 -181
rect 879 -147 945 -131
rect 879 -181 895 -147
rect 929 -181 945 -147
rect 879 -197 945 -181
rect 1071 -147 1137 -131
rect 1071 -181 1087 -147
rect 1121 -181 1137 -147
rect 1071 -197 1137 -181
rect 1263 -147 1329 -131
rect 1263 -181 1279 -147
rect 1313 -181 1329 -147
rect 1263 -197 1329 -181
<< polycont >>
rect -1313 147 -1279 181
rect -1121 147 -1087 181
rect -929 147 -895 181
rect -737 147 -703 181
rect -545 147 -511 181
rect -353 147 -319 181
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect 415 147 449 181
rect 607 147 641 181
rect 799 147 833 181
rect 991 147 1025 181
rect 1183 147 1217 181
rect 1375 147 1409 181
rect -1409 -181 -1375 -147
rect -1217 -181 -1183 -147
rect -1025 -181 -991 -147
rect -833 -181 -799 -147
rect -641 -181 -607 -147
rect -449 -181 -415 -147
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
rect 319 -181 353 -147
rect 511 -181 545 -147
rect 703 -181 737 -147
rect 895 -181 929 -147
rect 1087 -181 1121 -147
rect 1279 -181 1313 -147
<< locali >>
rect -1571 249 -1475 283
rect 1475 249 1571 283
rect -1571 187 -1537 249
rect 1537 187 1571 249
rect -1329 147 -1313 181
rect -1279 147 -1263 181
rect -1137 147 -1121 181
rect -1087 147 -1071 181
rect -945 147 -929 181
rect -895 147 -879 181
rect -753 147 -737 181
rect -703 147 -687 181
rect -561 147 -545 181
rect -511 147 -495 181
rect -369 147 -353 181
rect -319 147 -303 181
rect -177 147 -161 181
rect -127 147 -111 181
rect 15 147 31 181
rect 65 147 81 181
rect 207 147 223 181
rect 257 147 273 181
rect 399 147 415 181
rect 449 147 465 181
rect 591 147 607 181
rect 641 147 657 181
rect 783 147 799 181
rect 833 147 849 181
rect 975 147 991 181
rect 1025 147 1041 181
rect 1167 147 1183 181
rect 1217 147 1233 181
rect 1359 147 1375 181
rect 1409 147 1425 181
rect -1457 88 -1423 104
rect -1457 -104 -1423 -88
rect -1361 88 -1327 104
rect -1361 -104 -1327 -88
rect -1265 88 -1231 104
rect -1265 -104 -1231 -88
rect -1169 88 -1135 104
rect -1169 -104 -1135 -88
rect -1073 88 -1039 104
rect -1073 -104 -1039 -88
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -881 88 -847 104
rect -881 -104 -847 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -689 88 -655 104
rect -689 -104 -655 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 655 88 689 104
rect 655 -104 689 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 847 88 881 104
rect 847 -104 881 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect 1039 88 1073 104
rect 1039 -104 1073 -88
rect 1135 88 1169 104
rect 1135 -104 1169 -88
rect 1231 88 1265 104
rect 1231 -104 1265 -88
rect 1327 88 1361 104
rect 1327 -104 1361 -88
rect 1423 88 1457 104
rect 1423 -104 1457 -88
rect -1425 -181 -1409 -147
rect -1375 -181 -1359 -147
rect -1233 -181 -1217 -147
rect -1183 -181 -1167 -147
rect -1041 -181 -1025 -147
rect -991 -181 -975 -147
rect -849 -181 -833 -147
rect -799 -181 -783 -147
rect -657 -181 -641 -147
rect -607 -181 -591 -147
rect -465 -181 -449 -147
rect -415 -181 -399 -147
rect -273 -181 -257 -147
rect -223 -181 -207 -147
rect -81 -181 -65 -147
rect -31 -181 -15 -147
rect 111 -181 127 -147
rect 161 -181 177 -147
rect 303 -181 319 -147
rect 353 -181 369 -147
rect 495 -181 511 -147
rect 545 -181 561 -147
rect 687 -181 703 -147
rect 737 -181 753 -147
rect 879 -181 895 -147
rect 929 -181 945 -147
rect 1071 -181 1087 -147
rect 1121 -181 1137 -147
rect 1263 -181 1279 -147
rect 1313 -181 1329 -147
rect -1571 -249 -1537 -187
rect 1537 -249 1571 -187
rect -1571 -283 -1475 -249
rect 1475 -283 1571 -249
<< viali >>
rect -1313 147 -1279 181
rect -1121 147 -1087 181
rect -929 147 -895 181
rect -737 147 -703 181
rect -545 147 -511 181
rect -353 147 -319 181
rect -161 147 -127 181
rect 31 147 65 181
rect 223 147 257 181
rect 415 147 449 181
rect 607 147 641 181
rect 799 147 833 181
rect 991 147 1025 181
rect 1183 147 1217 181
rect 1375 147 1409 181
rect -1457 -88 -1423 88
rect -1361 -88 -1327 88
rect -1265 -88 -1231 88
rect -1169 -88 -1135 88
rect -1073 -88 -1039 88
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect 1039 -88 1073 88
rect 1135 -88 1169 88
rect 1231 -88 1265 88
rect 1327 -88 1361 88
rect 1423 -88 1457 88
rect -1409 -181 -1375 -147
rect -1217 -181 -1183 -147
rect -1025 -181 -991 -147
rect -833 -181 -799 -147
rect -641 -181 -607 -147
rect -449 -181 -415 -147
rect -257 -181 -223 -147
rect -65 -181 -31 -147
rect 127 -181 161 -147
rect 319 -181 353 -147
rect 511 -181 545 -147
rect 703 -181 737 -147
rect 895 -181 929 -147
rect 1087 -181 1121 -147
rect 1279 -181 1313 -147
<< metal1 >>
rect -1325 181 -1267 187
rect -1325 147 -1313 181
rect -1279 147 -1267 181
rect -1325 141 -1267 147
rect -1133 181 -1075 187
rect -1133 147 -1121 181
rect -1087 147 -1075 181
rect -1133 141 -1075 147
rect -941 181 -883 187
rect -941 147 -929 181
rect -895 147 -883 181
rect -941 141 -883 147
rect -749 181 -691 187
rect -749 147 -737 181
rect -703 147 -691 181
rect -749 141 -691 147
rect -557 181 -499 187
rect -557 147 -545 181
rect -511 147 -499 181
rect -557 141 -499 147
rect -365 181 -307 187
rect -365 147 -353 181
rect -319 147 -307 181
rect -365 141 -307 147
rect -173 181 -115 187
rect -173 147 -161 181
rect -127 147 -115 181
rect -173 141 -115 147
rect 19 181 77 187
rect 19 147 31 181
rect 65 147 77 181
rect 19 141 77 147
rect 211 181 269 187
rect 211 147 223 181
rect 257 147 269 181
rect 211 141 269 147
rect 403 181 461 187
rect 403 147 415 181
rect 449 147 461 181
rect 403 141 461 147
rect 595 181 653 187
rect 595 147 607 181
rect 641 147 653 181
rect 595 141 653 147
rect 787 181 845 187
rect 787 147 799 181
rect 833 147 845 181
rect 787 141 845 147
rect 979 181 1037 187
rect 979 147 991 181
rect 1025 147 1037 181
rect 979 141 1037 147
rect 1171 181 1229 187
rect 1171 147 1183 181
rect 1217 147 1229 181
rect 1171 141 1229 147
rect 1363 181 1421 187
rect 1363 147 1375 181
rect 1409 147 1421 181
rect 1363 141 1421 147
rect -1463 88 -1417 100
rect -1463 -88 -1457 88
rect -1423 -88 -1417 88
rect -1463 -100 -1417 -88
rect -1367 88 -1321 100
rect -1367 -88 -1361 88
rect -1327 -88 -1321 88
rect -1367 -100 -1321 -88
rect -1271 88 -1225 100
rect -1271 -88 -1265 88
rect -1231 -88 -1225 88
rect -1271 -100 -1225 -88
rect -1175 88 -1129 100
rect -1175 -88 -1169 88
rect -1135 -88 -1129 88
rect -1175 -100 -1129 -88
rect -1079 88 -1033 100
rect -1079 -88 -1073 88
rect -1039 -88 -1033 88
rect -1079 -100 -1033 -88
rect -983 88 -937 100
rect -983 -88 -977 88
rect -943 -88 -937 88
rect -983 -100 -937 -88
rect -887 88 -841 100
rect -887 -88 -881 88
rect -847 -88 -841 88
rect -887 -100 -841 -88
rect -791 88 -745 100
rect -791 -88 -785 88
rect -751 -88 -745 88
rect -791 -100 -745 -88
rect -695 88 -649 100
rect -695 -88 -689 88
rect -655 -88 -649 88
rect -695 -100 -649 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 649 88 695 100
rect 649 -88 655 88
rect 689 -88 695 88
rect 649 -100 695 -88
rect 745 88 791 100
rect 745 -88 751 88
rect 785 -88 791 88
rect 745 -100 791 -88
rect 841 88 887 100
rect 841 -88 847 88
rect 881 -88 887 88
rect 841 -100 887 -88
rect 937 88 983 100
rect 937 -88 943 88
rect 977 -88 983 88
rect 937 -100 983 -88
rect 1033 88 1079 100
rect 1033 -88 1039 88
rect 1073 -88 1079 88
rect 1033 -100 1079 -88
rect 1129 88 1175 100
rect 1129 -88 1135 88
rect 1169 -88 1175 88
rect 1129 -100 1175 -88
rect 1225 88 1271 100
rect 1225 -88 1231 88
rect 1265 -88 1271 88
rect 1225 -100 1271 -88
rect 1321 88 1367 100
rect 1321 -88 1327 88
rect 1361 -88 1367 88
rect 1321 -100 1367 -88
rect 1417 88 1463 100
rect 1417 -88 1423 88
rect 1457 -88 1463 88
rect 1417 -100 1463 -88
rect -1421 -147 -1363 -141
rect -1421 -181 -1409 -147
rect -1375 -181 -1363 -147
rect -1421 -187 -1363 -181
rect -1229 -147 -1171 -141
rect -1229 -181 -1217 -147
rect -1183 -181 -1171 -147
rect -1229 -187 -1171 -181
rect -1037 -147 -979 -141
rect -1037 -181 -1025 -147
rect -991 -181 -979 -147
rect -1037 -187 -979 -181
rect -845 -147 -787 -141
rect -845 -181 -833 -147
rect -799 -181 -787 -147
rect -845 -187 -787 -181
rect -653 -147 -595 -141
rect -653 -181 -641 -147
rect -607 -181 -595 -147
rect -653 -187 -595 -181
rect -461 -147 -403 -141
rect -461 -181 -449 -147
rect -415 -181 -403 -147
rect -461 -187 -403 -181
rect -269 -147 -211 -141
rect -269 -181 -257 -147
rect -223 -181 -211 -147
rect -269 -187 -211 -181
rect -77 -147 -19 -141
rect -77 -181 -65 -147
rect -31 -181 -19 -147
rect -77 -187 -19 -181
rect 115 -147 173 -141
rect 115 -181 127 -147
rect 161 -181 173 -147
rect 115 -187 173 -181
rect 307 -147 365 -141
rect 307 -181 319 -147
rect 353 -181 365 -147
rect 307 -187 365 -181
rect 499 -147 557 -141
rect 499 -181 511 -147
rect 545 -181 557 -147
rect 499 -187 557 -181
rect 691 -147 749 -141
rect 691 -181 703 -147
rect 737 -181 749 -147
rect 691 -187 749 -181
rect 883 -147 941 -141
rect 883 -181 895 -147
rect 929 -181 941 -147
rect 883 -187 941 -181
rect 1075 -147 1133 -141
rect 1075 -181 1087 -147
rect 1121 -181 1133 -147
rect 1075 -187 1133 -181
rect 1267 -147 1325 -141
rect 1267 -181 1279 -147
rect 1313 -181 1325 -147
rect 1267 -187 1325 -181
<< properties >>
string FIXED_BBOX -1554 -266 1554 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1 l 0.15 m 1 nf 30 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
