** sch_path: /home/ricardoatt/RATT_repos/Proyectos_xschem/opamp_design/folded_cascode_opamp/folded_one_stage_opamp_sr.sch
**.subckt folded_one_stage_opamp_sr
V1 VDD GND 1.8
V3 Vinp GND PWL(0 0 4.999u 0 5u 1.8 9.999u 1.8 10u 0)
V4 VSS GND 0
x1 VDD Vout Vinp Vout VSS folded_cascode_opamp
**** begin user architecture code


.param W1= 0.45
.param W3= 16.776
.param W4= 65.116
.param W8= 43.6
.param L0= 0.45
.control
	tran 0.1n 15u
	set color0=rgb:f/f/f
	set color1=rgb:0/0/0
	plot v(Vout)
	wrdata cascode_one_stage_opamp_sr.ssv (Vout)
.endc
.save all



.param mc_mm_switch=0
.param mc_pr_switch=0
.include /home/ricardoatt/pdk/sky130B/libs.tech/ngspice/corners/tt.spice
.include /home/ricardoatt/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical.spice
.include /home/ricardoatt/pdk/sky130B/libs.tech/ngspice/r+c/res_typical__cap_typical__lin.spice
.include /home/ricardoatt/pdk/sky130B/libs.tech/ngspice/corners/tt/specialized_cells.spice

**** end user architecture code
**.ends

* expanding   symbol:
*+  /home/ricardoatt/RATT_repos/Proyectos_xschem/opamp_design/folded_cascode_opamp/folded_cascode_opamp.sym # of pins=5
** sym_path: /home/ricardoatt/RATT_repos/Proyectos_xschem/opamp_design/folded_cascode_opamp/folded_cascode_opamp.sym
** sch_path: /home/ricardoatt/RATT_repos/Proyectos_xschem/opamp_design/folded_cascode_opamp/folded_cascode_opamp.sch
.subckt folded_cascode_opamp VDD Vout Vinp Vinn VSS
*.opin Vout
*.ipin Vinn
*.ipin Vinp
*.iopin VDD
*.iopin VSS
XM11 net4 net2 VSS VSS sky130_fd_pr__nfet_01v8 L={L0} W={W8} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 net3 net2 VSS VSS sky130_fd_pr__nfet_01v8 L={L0} W={W8} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net2 net1 net3 VSS sky130_fd_pr__nfet_01v8 L={L0} W={W8} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 Vout net1 net4 VSS sky130_fd_pr__nfet_01v8 L={L0} W={W8} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 Vout net5 net8 VDD sky130_fd_pr__pfet_01v8 L={L0} W={W4} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 net2 net5 net7 VDD sky130_fd_pr__pfet_01v8 L={L0} W={W4} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM1 net7 Vinp net6 VSS sky130_fd_pr__nfet_01v8 L={L0} W={W1} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net8 Vinn net6 VSS sky130_fd_pr__nfet_01v8 L={L0} W={W1} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net6 net10 VSS VSS sky130_fd_pr__nfet_01v8 L={L0} W={W3} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net7 net9 VDD VDD sky130_fd_pr__pfet_01v8 L={L0} W={W4} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net8 net9 VDD VDD sky130_fd_pr__pfet_01v8 L={L0} W={W4} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 net9 net9 VDD VDD sky130_fd_pr__pfet_01v8 L={L0} W={W4} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I4 net9 VSS 165u
XM13 net5 net5 VDD VDD sky130_fd_pr__pfet_01v8 L={L0} W={W4} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I1 net5 VSS 165u
XM14 net1 net1 VSS VSS sky130_fd_pr__nfet_01v8 L={L0} W={W8} nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
I2 VDD net1 165u
XM15 net10 net10 VSS VSS sky130_fd_pr__nfet_01v8 L={L0} W={W3} nf=1 ad='int((nf+1)/2) * W/nf * 0.29'
+ as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)'
+ nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
I3 VDD net10 150u
.ends

.GLOBAL VDD
.GLOBAL GND
.end
