magic
tech sky130B
magscale 1 2
timestamp 1727994832
<< error_p >>
rect -29 -511 29 -505
rect -29 -545 -17 -511
rect -29 -551 29 -545
<< nwell >>
rect -211 -684 211 684
<< pmos >>
rect -15 -464 15 536
<< pdiff >>
rect -73 524 -15 536
rect -73 -452 -61 524
rect -27 -452 -15 524
rect -73 -464 -15 -452
rect 15 524 73 536
rect 15 -452 27 524
rect 61 -452 73 524
rect 15 -464 73 -452
<< pdiffc >>
rect -61 -452 -27 524
rect 27 -452 61 524
<< nsubdiff >>
rect -175 614 -79 648
rect 79 614 175 648
rect -175 551 -141 614
rect 141 551 175 614
rect -175 -614 -141 -551
rect 141 -614 175 -551
rect -175 -648 -79 -614
rect 79 -648 175 -614
<< nsubdiffcont >>
rect -79 614 79 648
rect -175 -551 -141 551
rect 141 -551 175 551
rect -79 -648 79 -614
<< poly >>
rect -15 536 15 562
rect -15 -495 15 -464
rect -33 -511 33 -495
rect -33 -545 -17 -511
rect 17 -545 33 -511
rect -33 -561 33 -545
<< polycont >>
rect -17 -545 17 -511
<< locali >>
rect -175 614 -79 648
rect 79 614 175 648
rect -175 551 -141 614
rect 141 551 175 614
rect -61 524 -27 540
rect -61 -468 -27 -452
rect 27 524 61 540
rect 27 -468 61 -452
rect -33 -545 -17 -511
rect 17 -545 33 -511
rect -175 -614 -141 -551
rect 141 -614 175 -551
rect -175 -648 -79 -614
rect 79 -648 175 -614
<< viali >>
rect -61 -452 -27 524
rect 27 -452 61 524
rect -17 -545 17 -511
<< metal1 >>
rect -67 524 -21 536
rect -67 -452 -61 524
rect -27 -452 -21 524
rect -67 -464 -21 -452
rect 21 524 67 536
rect 21 -452 27 524
rect 61 -452 67 524
rect 21 -464 67 -452
rect -29 -511 29 -505
rect -29 -545 -17 -511
rect 17 -545 29 -511
rect -29 -551 29 -545
<< labels >>
flabel metal1 s 44 34 44 34 0 FreeSans 480 0 0 0 D
port 16 nsew
flabel metal1 s -44 36 -44 36 0 FreeSans 480 0 0 0 S
port 17 nsew
flabel metal1 s 0 -528 0 -528 0 FreeSans 480 0 0 0 G
port 18 nsew
flabel locali s 0 631 0 631 0 FreeSans 480 0 0 0 B
port 19 nsew
<< properties >>
string FIXED_BBOX -158 -631 158 631
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 5.0 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 0 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
