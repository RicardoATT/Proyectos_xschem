magic
tech sky130B
magscale 1 2
timestamp 1728345824
<< error_s >>
rect 298 1115 333 1132
rect 299 1114 333 1115
rect 299 1078 369 1114
rect 685 1078 738 1079
rect 129 1047 187 1053
rect 129 1013 141 1047
rect 316 1044 387 1078
rect 667 1044 738 1078
rect 129 1007 187 1013
rect 129 719 187 725
rect 129 685 141 719
rect 129 679 187 685
rect 316 583 386 1044
rect 668 1043 738 1044
rect 685 1009 756 1043
rect 1036 1009 1071 1026
rect 498 976 556 982
rect 498 942 510 976
rect 498 936 556 942
rect 498 666 556 672
rect 498 632 510 666
rect 498 626 556 632
rect 316 547 369 583
rect 685 530 755 1009
rect 1037 1008 1071 1009
rect 1037 972 1107 1008
rect 867 941 925 947
rect 867 907 879 941
rect 1054 938 1125 972
rect 1405 938 1440 972
rect 867 901 925 907
rect 867 613 925 619
rect 867 579 879 613
rect 867 573 925 579
rect 685 494 738 530
rect 1054 477 1124 938
rect 1406 919 1440 938
rect 1792 919 1845 920
rect 1236 870 1294 876
rect 1236 836 1248 870
rect 1236 830 1294 836
rect 1236 560 1294 566
rect 1236 526 1248 560
rect 1236 520 1294 526
rect 1054 441 1107 477
rect 1425 424 1440 919
rect 1459 885 1494 919
rect 1774 885 1845 919
rect 1459 424 1493 885
rect 1775 884 1845 885
rect 1792 850 1863 884
rect 2143 850 2178 884
rect 1605 817 1663 823
rect 1605 783 1617 817
rect 1605 777 1663 783
rect 1605 507 1663 513
rect 1605 473 1617 507
rect 1605 467 1663 473
rect 1459 390 1474 424
rect 1792 371 1862 850
rect 2144 831 2178 850
rect 1974 782 2032 788
rect 1974 748 1986 782
rect 1974 742 2032 748
rect 1974 454 2032 460
rect 1974 420 1986 454
rect 1974 414 2032 420
rect 1792 335 1845 371
rect 2163 318 2178 831
rect 2197 797 2232 831
rect 2512 797 2547 814
rect 2197 318 2231 797
rect 2513 796 2547 797
rect 2513 760 2583 796
rect 2899 760 2952 761
rect 2343 729 2401 735
rect 2343 695 2355 729
rect 2530 726 2601 760
rect 2881 726 2952 760
rect 2343 689 2401 695
rect 2343 401 2401 407
rect 2343 367 2355 401
rect 2343 361 2401 367
rect 2197 284 2212 318
rect 2530 265 2600 726
rect 2882 725 2952 726
rect 2899 691 2970 725
rect 3250 691 3285 725
rect 2712 658 2770 664
rect 2712 624 2724 658
rect 2712 618 2770 624
rect 2712 348 2770 354
rect 2712 314 2724 348
rect 2712 308 2770 314
rect 2530 229 2583 265
rect 2899 212 2969 691
rect 3251 672 3285 691
rect 3081 623 3139 629
rect 3081 589 3093 623
rect 3081 583 3139 589
rect 3081 295 3139 301
rect 3081 261 3093 295
rect 3081 255 3139 261
rect 2899 176 2952 212
rect 3270 159 3285 672
rect 3304 638 3339 672
rect 3619 638 3654 672
rect 3304 159 3338 638
rect 3620 619 3654 638
rect 3450 570 3508 576
rect 3450 536 3462 570
rect 3450 530 3508 536
rect 3450 242 3508 248
rect 3450 208 3462 242
rect 3450 202 3508 208
rect 3304 125 3319 159
rect 3639 106 3654 619
rect 3673 585 3708 619
rect 3988 585 4023 619
rect 3673 106 3707 585
rect 3989 566 4023 585
rect 3819 517 3877 523
rect 3819 483 3831 517
rect 3819 477 3877 483
rect 3819 189 3877 195
rect 3819 155 3831 189
rect 3819 149 3877 155
rect 3673 72 3688 106
rect 4008 53 4023 566
rect 4042 532 4077 566
rect 4357 532 4392 566
rect 4042 53 4076 532
rect 4358 513 4392 532
rect 4188 464 4246 470
rect 4188 430 4200 464
rect 4188 424 4246 430
rect 4188 136 4246 142
rect 4188 102 4200 136
rect 4188 96 4246 102
rect 4042 19 4057 53
rect 4377 0 4392 513
rect 4411 479 4446 513
rect 4726 479 4761 513
rect 4411 0 4445 479
rect 4727 460 4761 479
rect 4557 411 4615 417
rect 4557 377 4569 411
rect 4557 371 4615 377
rect 4557 83 4615 89
rect 4557 49 4569 83
rect 4557 43 4615 49
rect 4411 -34 4426 0
rect 4746 -53 4761 460
rect 4780 426 4815 460
rect 5095 426 5130 460
rect 4780 -53 4814 426
rect 5096 407 5130 426
rect 4926 358 4984 364
rect 4926 324 4938 358
rect 4926 318 4984 324
rect 4926 30 4984 36
rect 4926 -4 4938 30
rect 4926 -10 4984 -4
rect 4780 -87 4795 -53
rect 5115 -106 5130 407
rect 5149 373 5184 407
rect 5464 373 5499 390
rect 5149 -106 5183 373
rect 5465 372 5499 373
rect 5465 336 5535 372
rect 5295 305 5353 311
rect 5295 271 5307 305
rect 5482 302 5553 336
rect 5833 302 5868 336
rect 5295 265 5353 271
rect 5295 -23 5353 -17
rect 5295 -57 5307 -23
rect 5295 -63 5353 -57
rect 5149 -140 5164 -106
rect 5482 -159 5552 302
rect 5834 283 5868 302
rect 5664 234 5722 240
rect 5664 200 5676 234
rect 5664 194 5722 200
rect 5664 -76 5722 -70
rect 5664 -110 5676 -76
rect 5664 -116 5722 -110
rect 5482 -195 5535 -159
rect 5853 -212 5868 283
rect 5887 249 5922 283
rect 6202 249 6237 283
rect 5887 -212 5921 249
rect 6203 230 6237 249
rect 6033 181 6091 187
rect 6033 147 6045 181
rect 6033 141 6091 147
rect 6033 -129 6091 -123
rect 6033 -163 6045 -129
rect 6033 -169 6091 -163
rect 5887 -246 5902 -212
rect 6222 -265 6237 230
rect 6256 196 6291 230
rect 6571 196 6606 230
rect 6256 -265 6290 196
rect 6572 177 6606 196
rect 6402 128 6460 134
rect 6402 94 6414 128
rect 6402 88 6460 94
rect 6402 -182 6460 -176
rect 6402 -216 6414 -182
rect 6402 -222 6460 -216
rect 6256 -299 6271 -265
rect 6591 -318 6606 177
rect 6625 143 6660 177
rect 6940 143 6975 177
rect 6625 -318 6659 143
rect 6941 124 6975 143
rect 6771 75 6829 81
rect 6771 41 6783 75
rect 6771 35 6829 41
rect 6771 -235 6829 -229
rect 6771 -269 6783 -235
rect 6771 -275 6829 -269
rect 6625 -352 6640 -318
rect 6960 -371 6975 124
rect 6994 90 7029 124
rect 7309 90 7344 124
rect 6994 -371 7028 90
rect 7310 71 7344 90
rect 7140 22 7198 28
rect 7140 -12 7152 22
rect 7140 -18 7198 -12
rect 7140 -288 7198 -282
rect 7140 -322 7152 -288
rect 7140 -328 7198 -322
rect 6994 -405 7009 -371
rect 7329 -424 7344 71
rect 7363 37 7398 71
rect 7678 37 7713 71
rect 7363 -424 7397 37
rect 7679 18 7713 37
rect 8065 18 8118 19
rect 7509 -31 7567 -25
rect 7509 -65 7521 -31
rect 7509 -71 7567 -65
rect 7509 -341 7567 -335
rect 7509 -375 7521 -341
rect 7509 -381 7567 -375
rect 7363 -458 7378 -424
rect 7698 -477 7713 18
rect 7732 -16 7767 18
rect 8047 -16 8118 18
rect 7732 -477 7766 -16
rect 8048 -17 8118 -16
rect 8065 -51 8136 -17
rect 8416 -51 8451 -34
rect 7878 -84 7936 -78
rect 7878 -118 7890 -84
rect 7878 -124 7936 -118
rect 7878 -394 7936 -388
rect 7878 -428 7890 -394
rect 7878 -434 7936 -428
rect 7732 -511 7747 -477
rect 8065 -530 8135 -51
rect 8417 -52 8451 -51
rect 8417 -88 8487 -52
rect 8247 -119 8305 -113
rect 8247 -153 8259 -119
rect 8434 -122 8505 -88
rect 8247 -159 8305 -153
rect 8247 -447 8305 -441
rect 8247 -481 8259 -447
rect 8247 -487 8305 -481
rect 8065 -566 8118 -530
rect 8434 -583 8504 -122
rect 8616 -190 8674 -184
rect 8616 -224 8628 -190
rect 8616 -230 8674 -224
rect 8616 -500 8674 -494
rect 8616 -534 8628 -500
rect 8616 -540 8674 -534
rect 8434 -619 8487 -583
use sky130_fd_pr__pfet_01v8_XGS3BL  XM1
timestamp 1728345824
transform 1 0 2003 0 1 601
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1728345824
transform 1 0 1634 0 1 645
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM3
timestamp 1728345824
transform 1 0 896 0 1 760
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1728345824
transform 1 0 1265 0 1 698
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM5
timestamp 1728345824
transform 1 0 158 0 1 866
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM6
timestamp 1728345824
transform 1 0 527 0 1 804
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM7
timestamp 1728345824
transform 1 0 2372 0 1 548
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM8
timestamp 1728345824
transform 1 0 2741 0 1 486
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM9
timestamp 1728345824
transform 1 0 3110 0 1 442
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM10
timestamp 1728345824
transform 1 0 5693 0 1 62
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM11
timestamp 1728345824
transform 1 0 3479 0 1 389
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM12
timestamp 1728345824
transform 1 0 6062 0 1 9
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM13
timestamp 1728345824
transform 1 0 3848 0 1 336
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM14
timestamp 1728345824
transform 1 0 6431 0 1 -44
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM15
timestamp 1728345824
transform 1 0 4217 0 1 283
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM16
timestamp 1728345824
transform 1 0 6800 0 1 -97
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM17
timestamp 1728345824
transform 1 0 4586 0 1 230
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM18
timestamp 1728345824
transform 1 0 7169 0 1 -150
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM19
timestamp 1728345824
transform 1 0 4955 0 1 177
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM20
timestamp 1728345824
transform 1 0 7538 0 1 -203
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM21
timestamp 1728345824
transform 1 0 5324 0 1 124
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM22
timestamp 1728345824
transform 1 0 7907 0 1 -256
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM23
timestamp 1728345824
transform 1 0 8276 0 1 -300
box -211 -319 211 319
use sky130_fd_pr__nfet_01v8_648S5X  XM24
timestamp 1728345824
transform 1 0 8645 0 1 -362
box -211 -310 211 310
<< end >>
