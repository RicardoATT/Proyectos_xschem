magic
tech sky130B
magscale 1 2
timestamp 1729119800
<< error_p >>
rect -1085 201 -1027 207
rect -893 201 -835 207
rect -701 201 -643 207
rect -509 201 -451 207
rect -317 201 -259 207
rect -125 201 -67 207
rect 67 201 125 207
rect 259 201 317 207
rect 451 201 509 207
rect 643 201 701 207
rect 835 201 893 207
rect 1027 201 1085 207
rect -1085 167 -1073 201
rect -893 167 -881 201
rect -701 167 -689 201
rect -509 167 -497 201
rect -317 167 -305 201
rect -125 167 -113 201
rect 67 167 79 201
rect 259 167 271 201
rect 451 167 463 201
rect 643 167 655 201
rect 835 167 847 201
rect 1027 167 1039 201
rect -1085 161 -1027 167
rect -893 161 -835 167
rect -701 161 -643 167
rect -509 161 -451 167
rect -317 161 -259 167
rect -125 161 -67 167
rect 67 161 125 167
rect 259 161 317 167
rect 451 161 509 167
rect 643 161 701 167
rect 835 161 893 167
rect 1027 161 1085 167
rect -1181 -167 -1123 -161
rect -989 -167 -931 -161
rect -797 -167 -739 -161
rect -605 -167 -547 -161
rect -413 -167 -355 -161
rect -221 -167 -163 -161
rect -29 -167 29 -161
rect 163 -167 221 -161
rect 355 -167 413 -161
rect 547 -167 605 -161
rect 739 -167 797 -161
rect 931 -167 989 -161
rect 1123 -167 1181 -161
rect -1181 -201 -1169 -167
rect -989 -201 -977 -167
rect -797 -201 -785 -167
rect -605 -201 -593 -167
rect -413 -201 -401 -167
rect -221 -201 -209 -167
rect -29 -201 -17 -167
rect 163 -201 175 -167
rect 355 -201 367 -167
rect 547 -201 559 -167
rect 739 -201 751 -167
rect 931 -201 943 -167
rect 1123 -201 1135 -167
rect -1181 -207 -1123 -201
rect -989 -207 -931 -201
rect -797 -207 -739 -201
rect -605 -207 -547 -201
rect -413 -207 -355 -201
rect -221 -207 -163 -201
rect -29 -207 29 -201
rect 163 -207 221 -201
rect 355 -207 413 -201
rect 547 -207 605 -201
rect 739 -207 797 -201
rect 931 -207 989 -201
rect 1123 -207 1181 -201
<< nwell >>
rect -1367 -339 1367 339
<< pmos >>
rect -1167 -120 -1137 120
rect -1071 -120 -1041 120
rect -975 -120 -945 120
rect -879 -120 -849 120
rect -783 -120 -753 120
rect -687 -120 -657 120
rect -591 -120 -561 120
rect -495 -120 -465 120
rect -399 -120 -369 120
rect -303 -120 -273 120
rect -207 -120 -177 120
rect -111 -120 -81 120
rect -15 -120 15 120
rect 81 -120 111 120
rect 177 -120 207 120
rect 273 -120 303 120
rect 369 -120 399 120
rect 465 -120 495 120
rect 561 -120 591 120
rect 657 -120 687 120
rect 753 -120 783 120
rect 849 -120 879 120
rect 945 -120 975 120
rect 1041 -120 1071 120
rect 1137 -120 1167 120
<< pdiff >>
rect -1229 108 -1167 120
rect -1229 -108 -1217 108
rect -1183 -108 -1167 108
rect -1229 -120 -1167 -108
rect -1137 108 -1071 120
rect -1137 -108 -1121 108
rect -1087 -108 -1071 108
rect -1137 -120 -1071 -108
rect -1041 108 -975 120
rect -1041 -108 -1025 108
rect -991 -108 -975 108
rect -1041 -120 -975 -108
rect -945 108 -879 120
rect -945 -108 -929 108
rect -895 -108 -879 108
rect -945 -120 -879 -108
rect -849 108 -783 120
rect -849 -108 -833 108
rect -799 -108 -783 108
rect -849 -120 -783 -108
rect -753 108 -687 120
rect -753 -108 -737 108
rect -703 -108 -687 108
rect -753 -120 -687 -108
rect -657 108 -591 120
rect -657 -108 -641 108
rect -607 -108 -591 108
rect -657 -120 -591 -108
rect -561 108 -495 120
rect -561 -108 -545 108
rect -511 -108 -495 108
rect -561 -120 -495 -108
rect -465 108 -399 120
rect -465 -108 -449 108
rect -415 -108 -399 108
rect -465 -120 -399 -108
rect -369 108 -303 120
rect -369 -108 -353 108
rect -319 -108 -303 108
rect -369 -120 -303 -108
rect -273 108 -207 120
rect -273 -108 -257 108
rect -223 -108 -207 108
rect -273 -120 -207 -108
rect -177 108 -111 120
rect -177 -108 -161 108
rect -127 -108 -111 108
rect -177 -120 -111 -108
rect -81 108 -15 120
rect -81 -108 -65 108
rect -31 -108 -15 108
rect -81 -120 -15 -108
rect 15 108 81 120
rect 15 -108 31 108
rect 65 -108 81 108
rect 15 -120 81 -108
rect 111 108 177 120
rect 111 -108 127 108
rect 161 -108 177 108
rect 111 -120 177 -108
rect 207 108 273 120
rect 207 -108 223 108
rect 257 -108 273 108
rect 207 -120 273 -108
rect 303 108 369 120
rect 303 -108 319 108
rect 353 -108 369 108
rect 303 -120 369 -108
rect 399 108 465 120
rect 399 -108 415 108
rect 449 -108 465 108
rect 399 -120 465 -108
rect 495 108 561 120
rect 495 -108 511 108
rect 545 -108 561 108
rect 495 -120 561 -108
rect 591 108 657 120
rect 591 -108 607 108
rect 641 -108 657 108
rect 591 -120 657 -108
rect 687 108 753 120
rect 687 -108 703 108
rect 737 -108 753 108
rect 687 -120 753 -108
rect 783 108 849 120
rect 783 -108 799 108
rect 833 -108 849 108
rect 783 -120 849 -108
rect 879 108 945 120
rect 879 -108 895 108
rect 929 -108 945 108
rect 879 -120 945 -108
rect 975 108 1041 120
rect 975 -108 991 108
rect 1025 -108 1041 108
rect 975 -120 1041 -108
rect 1071 108 1137 120
rect 1071 -108 1087 108
rect 1121 -108 1137 108
rect 1071 -120 1137 -108
rect 1167 108 1229 120
rect 1167 -108 1183 108
rect 1217 -108 1229 108
rect 1167 -120 1229 -108
<< pdiffc >>
rect -1217 -108 -1183 108
rect -1121 -108 -1087 108
rect -1025 -108 -991 108
rect -929 -108 -895 108
rect -833 -108 -799 108
rect -737 -108 -703 108
rect -641 -108 -607 108
rect -545 -108 -511 108
rect -449 -108 -415 108
rect -353 -108 -319 108
rect -257 -108 -223 108
rect -161 -108 -127 108
rect -65 -108 -31 108
rect 31 -108 65 108
rect 127 -108 161 108
rect 223 -108 257 108
rect 319 -108 353 108
rect 415 -108 449 108
rect 511 -108 545 108
rect 607 -108 641 108
rect 703 -108 737 108
rect 799 -108 833 108
rect 895 -108 929 108
rect 991 -108 1025 108
rect 1087 -108 1121 108
rect 1183 -108 1217 108
<< nsubdiff >>
rect -1331 269 -1235 303
rect 1235 269 1331 303
rect -1331 207 -1297 269
rect 1297 207 1331 269
rect -1331 -269 -1297 -207
rect 1297 -269 1331 -207
rect -1331 -303 -1235 -269
rect 1235 -303 1331 -269
<< nsubdiffcont >>
rect -1235 269 1235 303
rect -1331 -207 -1297 207
rect 1297 -207 1331 207
rect -1235 -303 1235 -269
<< poly >>
rect -1089 201 -1023 217
rect -1089 167 -1073 201
rect -1039 167 -1023 201
rect -1089 151 -1023 167
rect -897 201 -831 217
rect -897 167 -881 201
rect -847 167 -831 201
rect -897 151 -831 167
rect -705 201 -639 217
rect -705 167 -689 201
rect -655 167 -639 201
rect -705 151 -639 167
rect -513 201 -447 217
rect -513 167 -497 201
rect -463 167 -447 201
rect -513 151 -447 167
rect -321 201 -255 217
rect -321 167 -305 201
rect -271 167 -255 201
rect -321 151 -255 167
rect -129 201 -63 217
rect -129 167 -113 201
rect -79 167 -63 201
rect -129 151 -63 167
rect 63 201 129 217
rect 63 167 79 201
rect 113 167 129 201
rect 63 151 129 167
rect 255 201 321 217
rect 255 167 271 201
rect 305 167 321 201
rect 255 151 321 167
rect 447 201 513 217
rect 447 167 463 201
rect 497 167 513 201
rect 447 151 513 167
rect 639 201 705 217
rect 639 167 655 201
rect 689 167 705 201
rect 639 151 705 167
rect 831 201 897 217
rect 831 167 847 201
rect 881 167 897 201
rect 831 151 897 167
rect 1023 201 1089 217
rect 1023 167 1039 201
rect 1073 167 1089 201
rect 1023 151 1089 167
rect -1167 120 -1137 146
rect -1071 120 -1041 151
rect -975 120 -945 146
rect -879 120 -849 151
rect -783 120 -753 146
rect -687 120 -657 151
rect -591 120 -561 146
rect -495 120 -465 151
rect -399 120 -369 146
rect -303 120 -273 151
rect -207 120 -177 146
rect -111 120 -81 151
rect -15 120 15 146
rect 81 120 111 151
rect 177 120 207 146
rect 273 120 303 151
rect 369 120 399 146
rect 465 120 495 151
rect 561 120 591 146
rect 657 120 687 151
rect 753 120 783 146
rect 849 120 879 151
rect 945 120 975 146
rect 1041 120 1071 151
rect 1137 120 1167 146
rect -1167 -151 -1137 -120
rect -1071 -146 -1041 -120
rect -975 -151 -945 -120
rect -879 -146 -849 -120
rect -783 -151 -753 -120
rect -687 -146 -657 -120
rect -591 -151 -561 -120
rect -495 -146 -465 -120
rect -399 -151 -369 -120
rect -303 -146 -273 -120
rect -207 -151 -177 -120
rect -111 -146 -81 -120
rect -15 -151 15 -120
rect 81 -146 111 -120
rect 177 -151 207 -120
rect 273 -146 303 -120
rect 369 -151 399 -120
rect 465 -146 495 -120
rect 561 -151 591 -120
rect 657 -146 687 -120
rect 753 -151 783 -120
rect 849 -146 879 -120
rect 945 -151 975 -120
rect 1041 -146 1071 -120
rect 1137 -151 1167 -120
rect -1185 -167 -1119 -151
rect -1185 -201 -1169 -167
rect -1135 -201 -1119 -167
rect -1185 -217 -1119 -201
rect -993 -167 -927 -151
rect -993 -201 -977 -167
rect -943 -201 -927 -167
rect -993 -217 -927 -201
rect -801 -167 -735 -151
rect -801 -201 -785 -167
rect -751 -201 -735 -167
rect -801 -217 -735 -201
rect -609 -167 -543 -151
rect -609 -201 -593 -167
rect -559 -201 -543 -167
rect -609 -217 -543 -201
rect -417 -167 -351 -151
rect -417 -201 -401 -167
rect -367 -201 -351 -167
rect -417 -217 -351 -201
rect -225 -167 -159 -151
rect -225 -201 -209 -167
rect -175 -201 -159 -167
rect -225 -217 -159 -201
rect -33 -167 33 -151
rect -33 -201 -17 -167
rect 17 -201 33 -167
rect -33 -217 33 -201
rect 159 -167 225 -151
rect 159 -201 175 -167
rect 209 -201 225 -167
rect 159 -217 225 -201
rect 351 -167 417 -151
rect 351 -201 367 -167
rect 401 -201 417 -167
rect 351 -217 417 -201
rect 543 -167 609 -151
rect 543 -201 559 -167
rect 593 -201 609 -167
rect 543 -217 609 -201
rect 735 -167 801 -151
rect 735 -201 751 -167
rect 785 -201 801 -167
rect 735 -217 801 -201
rect 927 -167 993 -151
rect 927 -201 943 -167
rect 977 -201 993 -167
rect 927 -217 993 -201
rect 1119 -167 1185 -151
rect 1119 -201 1135 -167
rect 1169 -201 1185 -167
rect 1119 -217 1185 -201
<< polycont >>
rect -1073 167 -1039 201
rect -881 167 -847 201
rect -689 167 -655 201
rect -497 167 -463 201
rect -305 167 -271 201
rect -113 167 -79 201
rect 79 167 113 201
rect 271 167 305 201
rect 463 167 497 201
rect 655 167 689 201
rect 847 167 881 201
rect 1039 167 1073 201
rect -1169 -201 -1135 -167
rect -977 -201 -943 -167
rect -785 -201 -751 -167
rect -593 -201 -559 -167
rect -401 -201 -367 -167
rect -209 -201 -175 -167
rect -17 -201 17 -167
rect 175 -201 209 -167
rect 367 -201 401 -167
rect 559 -201 593 -167
rect 751 -201 785 -167
rect 943 -201 977 -167
rect 1135 -201 1169 -167
<< locali >>
rect -1331 269 -1235 303
rect 1235 269 1331 303
rect -1331 207 -1297 269
rect 1297 207 1331 269
rect -1089 167 -1073 201
rect -1039 167 -1023 201
rect -897 167 -881 201
rect -847 167 -831 201
rect -705 167 -689 201
rect -655 167 -639 201
rect -513 167 -497 201
rect -463 167 -447 201
rect -321 167 -305 201
rect -271 167 -255 201
rect -129 167 -113 201
rect -79 167 -63 201
rect 63 167 79 201
rect 113 167 129 201
rect 255 167 271 201
rect 305 167 321 201
rect 447 167 463 201
rect 497 167 513 201
rect 639 167 655 201
rect 689 167 705 201
rect 831 167 847 201
rect 881 167 897 201
rect 1023 167 1039 201
rect 1073 167 1089 201
rect -1217 108 -1183 124
rect -1217 -124 -1183 -108
rect -1121 108 -1087 124
rect -1121 -124 -1087 -108
rect -1025 108 -991 124
rect -1025 -124 -991 -108
rect -929 108 -895 124
rect -929 -124 -895 -108
rect -833 108 -799 124
rect -833 -124 -799 -108
rect -737 108 -703 124
rect -737 -124 -703 -108
rect -641 108 -607 124
rect -641 -124 -607 -108
rect -545 108 -511 124
rect -545 -124 -511 -108
rect -449 108 -415 124
rect -449 -124 -415 -108
rect -353 108 -319 124
rect -353 -124 -319 -108
rect -257 108 -223 124
rect -257 -124 -223 -108
rect -161 108 -127 124
rect -161 -124 -127 -108
rect -65 108 -31 124
rect -65 -124 -31 -108
rect 31 108 65 124
rect 31 -124 65 -108
rect 127 108 161 124
rect 127 -124 161 -108
rect 223 108 257 124
rect 223 -124 257 -108
rect 319 108 353 124
rect 319 -124 353 -108
rect 415 108 449 124
rect 415 -124 449 -108
rect 511 108 545 124
rect 511 -124 545 -108
rect 607 108 641 124
rect 607 -124 641 -108
rect 703 108 737 124
rect 703 -124 737 -108
rect 799 108 833 124
rect 799 -124 833 -108
rect 895 108 929 124
rect 895 -124 929 -108
rect 991 108 1025 124
rect 991 -124 1025 -108
rect 1087 108 1121 124
rect 1087 -124 1121 -108
rect 1183 108 1217 124
rect 1183 -124 1217 -108
rect -1185 -201 -1169 -167
rect -1135 -201 -1119 -167
rect -993 -201 -977 -167
rect -943 -201 -927 -167
rect -801 -201 -785 -167
rect -751 -201 -735 -167
rect -609 -201 -593 -167
rect -559 -201 -543 -167
rect -417 -201 -401 -167
rect -367 -201 -351 -167
rect -225 -201 -209 -167
rect -175 -201 -159 -167
rect -33 -201 -17 -167
rect 17 -201 33 -167
rect 159 -201 175 -167
rect 209 -201 225 -167
rect 351 -201 367 -167
rect 401 -201 417 -167
rect 543 -201 559 -167
rect 593 -201 609 -167
rect 735 -201 751 -167
rect 785 -201 801 -167
rect 927 -201 943 -167
rect 977 -201 993 -167
rect 1119 -201 1135 -167
rect 1169 -201 1185 -167
rect -1331 -269 -1297 -207
rect 1297 -269 1331 -207
rect -1331 -303 -1235 -269
rect 1235 -303 1331 -269
<< viali >>
rect -1073 167 -1039 201
rect -881 167 -847 201
rect -689 167 -655 201
rect -497 167 -463 201
rect -305 167 -271 201
rect -113 167 -79 201
rect 79 167 113 201
rect 271 167 305 201
rect 463 167 497 201
rect 655 167 689 201
rect 847 167 881 201
rect 1039 167 1073 201
rect -1217 -108 -1183 108
rect -1121 -108 -1087 108
rect -1025 -108 -991 108
rect -929 -108 -895 108
rect -833 -108 -799 108
rect -737 -108 -703 108
rect -641 -108 -607 108
rect -545 -108 -511 108
rect -449 -108 -415 108
rect -353 -108 -319 108
rect -257 -108 -223 108
rect -161 -108 -127 108
rect -65 -108 -31 108
rect 31 -108 65 108
rect 127 -108 161 108
rect 223 -108 257 108
rect 319 -108 353 108
rect 415 -108 449 108
rect 511 -108 545 108
rect 607 -108 641 108
rect 703 -108 737 108
rect 799 -108 833 108
rect 895 -108 929 108
rect 991 -108 1025 108
rect 1087 -108 1121 108
rect 1183 -108 1217 108
rect -1169 -201 -1135 -167
rect -977 -201 -943 -167
rect -785 -201 -751 -167
rect -593 -201 -559 -167
rect -401 -201 -367 -167
rect -209 -201 -175 -167
rect -17 -201 17 -167
rect 175 -201 209 -167
rect 367 -201 401 -167
rect 559 -201 593 -167
rect 751 -201 785 -167
rect 943 -201 977 -167
rect 1135 -201 1169 -167
<< metal1 >>
rect -1085 201 -1027 207
rect -1085 167 -1073 201
rect -1039 167 -1027 201
rect -1085 161 -1027 167
rect -893 201 -835 207
rect -893 167 -881 201
rect -847 167 -835 201
rect -893 161 -835 167
rect -701 201 -643 207
rect -701 167 -689 201
rect -655 167 -643 201
rect -701 161 -643 167
rect -509 201 -451 207
rect -509 167 -497 201
rect -463 167 -451 201
rect -509 161 -451 167
rect -317 201 -259 207
rect -317 167 -305 201
rect -271 167 -259 201
rect -317 161 -259 167
rect -125 201 -67 207
rect -125 167 -113 201
rect -79 167 -67 201
rect -125 161 -67 167
rect 67 201 125 207
rect 67 167 79 201
rect 113 167 125 201
rect 67 161 125 167
rect 259 201 317 207
rect 259 167 271 201
rect 305 167 317 201
rect 259 161 317 167
rect 451 201 509 207
rect 451 167 463 201
rect 497 167 509 201
rect 451 161 509 167
rect 643 201 701 207
rect 643 167 655 201
rect 689 167 701 201
rect 643 161 701 167
rect 835 201 893 207
rect 835 167 847 201
rect 881 167 893 201
rect 835 161 893 167
rect 1027 201 1085 207
rect 1027 167 1039 201
rect 1073 167 1085 201
rect 1027 161 1085 167
rect -1223 108 -1177 120
rect -1223 -108 -1217 108
rect -1183 -108 -1177 108
rect -1223 -120 -1177 -108
rect -1127 108 -1081 120
rect -1127 -108 -1121 108
rect -1087 -108 -1081 108
rect -1127 -120 -1081 -108
rect -1031 108 -985 120
rect -1031 -108 -1025 108
rect -991 -108 -985 108
rect -1031 -120 -985 -108
rect -935 108 -889 120
rect -935 -108 -929 108
rect -895 -108 -889 108
rect -935 -120 -889 -108
rect -839 108 -793 120
rect -839 -108 -833 108
rect -799 -108 -793 108
rect -839 -120 -793 -108
rect -743 108 -697 120
rect -743 -108 -737 108
rect -703 -108 -697 108
rect -743 -120 -697 -108
rect -647 108 -601 120
rect -647 -108 -641 108
rect -607 -108 -601 108
rect -647 -120 -601 -108
rect -551 108 -505 120
rect -551 -108 -545 108
rect -511 -108 -505 108
rect -551 -120 -505 -108
rect -455 108 -409 120
rect -455 -108 -449 108
rect -415 -108 -409 108
rect -455 -120 -409 -108
rect -359 108 -313 120
rect -359 -108 -353 108
rect -319 -108 -313 108
rect -359 -120 -313 -108
rect -263 108 -217 120
rect -263 -108 -257 108
rect -223 -108 -217 108
rect -263 -120 -217 -108
rect -167 108 -121 120
rect -167 -108 -161 108
rect -127 -108 -121 108
rect -167 -120 -121 -108
rect -71 108 -25 120
rect -71 -108 -65 108
rect -31 -108 -25 108
rect -71 -120 -25 -108
rect 25 108 71 120
rect 25 -108 31 108
rect 65 -108 71 108
rect 25 -120 71 -108
rect 121 108 167 120
rect 121 -108 127 108
rect 161 -108 167 108
rect 121 -120 167 -108
rect 217 108 263 120
rect 217 -108 223 108
rect 257 -108 263 108
rect 217 -120 263 -108
rect 313 108 359 120
rect 313 -108 319 108
rect 353 -108 359 108
rect 313 -120 359 -108
rect 409 108 455 120
rect 409 -108 415 108
rect 449 -108 455 108
rect 409 -120 455 -108
rect 505 108 551 120
rect 505 -108 511 108
rect 545 -108 551 108
rect 505 -120 551 -108
rect 601 108 647 120
rect 601 -108 607 108
rect 641 -108 647 108
rect 601 -120 647 -108
rect 697 108 743 120
rect 697 -108 703 108
rect 737 -108 743 108
rect 697 -120 743 -108
rect 793 108 839 120
rect 793 -108 799 108
rect 833 -108 839 108
rect 793 -120 839 -108
rect 889 108 935 120
rect 889 -108 895 108
rect 929 -108 935 108
rect 889 -120 935 -108
rect 985 108 1031 120
rect 985 -108 991 108
rect 1025 -108 1031 108
rect 985 -120 1031 -108
rect 1081 108 1127 120
rect 1081 -108 1087 108
rect 1121 -108 1127 108
rect 1081 -120 1127 -108
rect 1177 108 1223 120
rect 1177 -108 1183 108
rect 1217 -108 1223 108
rect 1177 -120 1223 -108
rect -1181 -167 -1123 -161
rect -1181 -201 -1169 -167
rect -1135 -201 -1123 -167
rect -1181 -207 -1123 -201
rect -989 -167 -931 -161
rect -989 -201 -977 -167
rect -943 -201 -931 -167
rect -989 -207 -931 -201
rect -797 -167 -739 -161
rect -797 -201 -785 -167
rect -751 -201 -739 -167
rect -797 -207 -739 -201
rect -605 -167 -547 -161
rect -605 -201 -593 -167
rect -559 -201 -547 -167
rect -605 -207 -547 -201
rect -413 -167 -355 -161
rect -413 -201 -401 -167
rect -367 -201 -355 -167
rect -413 -207 -355 -201
rect -221 -167 -163 -161
rect -221 -201 -209 -167
rect -175 -201 -163 -167
rect -221 -207 -163 -201
rect -29 -167 29 -161
rect -29 -201 -17 -167
rect 17 -201 29 -167
rect -29 -207 29 -201
rect 163 -167 221 -161
rect 163 -201 175 -167
rect 209 -201 221 -167
rect 163 -207 221 -201
rect 355 -167 413 -161
rect 355 -201 367 -167
rect 401 -201 413 -167
rect 355 -207 413 -201
rect 547 -167 605 -161
rect 547 -201 559 -167
rect 593 -201 605 -167
rect 547 -207 605 -201
rect 739 -167 797 -161
rect 739 -201 751 -167
rect 785 -201 797 -167
rect 739 -207 797 -201
rect 931 -167 989 -161
rect 931 -201 943 -167
rect 977 -201 989 -167
rect 931 -207 989 -201
rect 1123 -167 1181 -161
rect 1123 -201 1135 -167
rect 1169 -201 1181 -167
rect 1123 -207 1181 -201
<< labels >>
flabel metal1 s -1056 184 -1056 184 0 FreeSans 480 0 0 0 G
port 8 nsew
flabel metal1 s -1200 1 -1200 1 0 FreeSans 480 0 0 0 D
port 9 nsew
flabel metal1 s -1103 -1 -1103 -1 0 FreeSans 480 0 0 0 S
port 10 nsew
flabel locali s -1 286 -1 286 0 FreeSans 480 0 0 0 B
port 11 nsew
<< properties >>
string FIXED_BBOX -1314 -286 1314 286
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.2 l 0.15 m 1 nf 25 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
